module DFC_TableA(
  input         clock,
  input         reset,
  output        io_cpu_w_data_ready,
  input         io_cpu_w_data_valid,
  input  [31:0] io_cpu_w_data_bits_listenAddr,
  input  [15:0] io_cpu_w_data_bits_wPid,
  output        io_cpu_l_data_ready,
  input         io_cpu_l_data_valid,
  input  [31:0] io_cpu_l_data_bits_listenAddr,
  input         io_tableD_wdata_ready,
  output        io_tableD_wdata_valid,
  output [31:0] io_tableD_wdata_bits_listenAddr,
  output [5:0]  io_tableD_wdata_bits_tableAId,
  input         io_tableD_ldata_ready,
  output        io_tableD_ldata_valid,
  output [31:0] io_tableD_ldata_bits_listenAddr,
  output        io_tableD_wresp_ready,
  input         io_tableD_wresp_valid,
  input         io_tableD_wresp_bits,
  output        io_tableD_lresp_ready,
  input         io_tableD_lresp_valid,
  input  [5:0]  io_tableD_lresp_bits_tableAId,
  input         io_tableD_lresp_bits_finish,
  input         io_cpu_expt_data_ready,
  output        io_cpu_expt_data_valid,
  output [15:0] io_cpu_expt_data_bits_pid,
  output        io_dfc_full_data_valid,
  output        io_dfc_full_data_bits_full_sig
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] infoMetaMem_pid [0:63]; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_1_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_1_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_2_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_2_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_3_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_3_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_4_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_4_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_5_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_5_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_6_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_6_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_7_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_7_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_8_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_8_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_9_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_9_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_10_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_10_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_11_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_11_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_12_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_12_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_13_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_13_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_14_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_14_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_15_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_15_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_16_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_16_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_17_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_17_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_18_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_18_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_19_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_19_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_20_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_20_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_21_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_21_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_22_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_22_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_23_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_23_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_24_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_24_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_25_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_25_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_26_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_26_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_27_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_27_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_28_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_28_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_29_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_29_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_30_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_30_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_31_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_31_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_32_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_32_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_33_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_33_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_34_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_34_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_35_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_35_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_36_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_36_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_37_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_37_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_38_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_38_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_39_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_39_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_40_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_40_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_41_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_41_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_42_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_42_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_43_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_43_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_44_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_44_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_45_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_45_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_46_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_46_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_47_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_47_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_48_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_48_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_49_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_49_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_50_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_50_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_51_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_51_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_52_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_52_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_53_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_53_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_54_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_54_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_55_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_55_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_56_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_56_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_57_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_57_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_58_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_58_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_59_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_59_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_60_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_60_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_61_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_61_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_62_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_62_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_64_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_64_addr; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_63_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_63_addr; // @[DFCTableA.scala 30:32]
  wire  infoMetaMem_pid_MPORT_63_mask; // @[DFCTableA.scala 30:32]
  wire  infoMetaMem_pid_MPORT_63_en; // @[DFCTableA.scala 30:32]
  wire [15:0] infoMetaMem_pid_MPORT_65_data; // @[DFCTableA.scala 30:32]
  wire [5:0] infoMetaMem_pid_MPORT_65_addr; // @[DFCTableA.scala 30:32]
  wire  infoMetaMem_pid_MPORT_65_mask; // @[DFCTableA.scala 30:32]
  wire  infoMetaMem_pid_MPORT_65_en; // @[DFCTableA.scala 30:32]
  reg  infoMetaMem_pid_MPORT_64_en_pipe_0;
  reg [5:0] infoMetaMem_pid_MPORT_64_addr_pipe_0;
  reg [7:0] counter_0; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_1; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_2; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_3; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_4; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_5; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_6; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_7; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_8; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_9; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_10; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_11; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_12; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_13; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_14; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_15; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_16; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_17; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_18; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_19; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_20; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_21; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_22; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_23; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_24; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_25; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_26; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_27; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_28; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_29; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_30; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_31; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_32; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_33; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_34; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_35; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_36; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_37; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_38; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_39; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_40; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_41; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_42; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_43; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_44; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_45; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_46; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_47; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_48; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_49; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_50; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_51; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_52; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_53; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_54; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_55; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_56; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_57; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_58; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_59; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_60; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_61; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_62; // @[DFCTableA.scala 29:20]
  reg [7:0] counter_63; // @[DFCTableA.scala 29:20]
  reg [63:0] tableA_valid; // @[DFCTableA.scala 31:29]
  reg [3:0] state; // @[DFCTableA.scala 34:22]
  reg [3:0] laststate; // @[DFCTableA.scala 35:26]
  wire  is_idle = state == 4'h0; // @[DFCTableA.scala 36:23]
  reg [31:0] laddr_reg; // @[DFCTableA.scala 39:26]
  reg [15:0] pid_reg; // @[DFCTableA.scala 40:24]
  reg [15:0] pid_act; // @[DFCTableA.scala 41:24]
  reg [5:0] table_wId; // @[DFCTableA.scala 42:26]
  reg  full_a; // @[DFCTableA.scala 43:23]
  reg  full_a_last; // @[DFCTableA.scala 44:28]
  reg  full_d; // @[DFCTableA.scala 45:23]
  reg  full_d_last; // @[DFCTableA.scala 46:28]
  wire  wEn = is_idle & io_cpu_w_data_valid; // @[DFCTableA.scala 48:21]
  wire  _T_13 = ~full_a_last & ~full_d_last; // @[DFCTableA.scala 67:44]
  wire  _T_14 = full_a | full_d; // @[DFCTableA.scala 67:72]
  wire  _T_15 = ~full_a_last & ~full_d_last & (full_a | full_d); // @[DFCTableA.scala 67:61]
  wire  _T_23 = tableA_valid[1] ? 1'h0 : 1'h1; // @[DFCTableA.scala 79:21]
  wire [1:0] _T_25 = tableA_valid[2] ? {{1'd0}, _T_23} : 2'h2; // @[DFCTableA.scala 79:21]
  wire [1:0] _T_27 = tableA_valid[3] ? _T_25 : 2'h3; // @[DFCTableA.scala 79:21]
  wire [2:0] _T_29 = tableA_valid[4] ? {{1'd0}, _T_27} : 3'h4; // @[DFCTableA.scala 79:21]
  wire [2:0] _T_31 = tableA_valid[5] ? _T_29 : 3'h5; // @[DFCTableA.scala 79:21]
  wire [2:0] _T_33 = tableA_valid[6] ? _T_31 : 3'h6; // @[DFCTableA.scala 79:21]
  wire [2:0] _T_35 = tableA_valid[7] ? _T_33 : 3'h7; // @[DFCTableA.scala 79:21]
  wire [3:0] _T_37 = tableA_valid[8] ? {{1'd0}, _T_35} : 4'h8; // @[DFCTableA.scala 79:21]
  wire [3:0] _T_39 = tableA_valid[9] ? _T_37 : 4'h9; // @[DFCTableA.scala 79:21]
  wire [3:0] _T_41 = tableA_valid[10] ? _T_39 : 4'ha; // @[DFCTableA.scala 79:21]
  wire [3:0] _T_43 = tableA_valid[11] ? _T_41 : 4'hb; // @[DFCTableA.scala 79:21]
  wire [3:0] _T_45 = tableA_valid[12] ? _T_43 : 4'hc; // @[DFCTableA.scala 79:21]
  wire [3:0] _T_47 = tableA_valid[13] ? _T_45 : 4'hd; // @[DFCTableA.scala 79:21]
  wire [3:0] _T_49 = tableA_valid[14] ? _T_47 : 4'he; // @[DFCTableA.scala 79:21]
  wire [3:0] _T_51 = tableA_valid[15] ? _T_49 : 4'hf; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_53 = tableA_valid[16] ? {{1'd0}, _T_51} : 5'h10; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_55 = tableA_valid[17] ? _T_53 : 5'h11; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_57 = tableA_valid[18] ? _T_55 : 5'h12; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_59 = tableA_valid[19] ? _T_57 : 5'h13; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_61 = tableA_valid[20] ? _T_59 : 5'h14; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_63 = tableA_valid[21] ? _T_61 : 5'h15; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_65 = tableA_valid[22] ? _T_63 : 5'h16; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_67 = tableA_valid[23] ? _T_65 : 5'h17; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_69 = tableA_valid[24] ? _T_67 : 5'h18; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_71 = tableA_valid[25] ? _T_69 : 5'h19; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_73 = tableA_valid[26] ? _T_71 : 5'h1a; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_75 = tableA_valid[27] ? _T_73 : 5'h1b; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_77 = tableA_valid[28] ? _T_75 : 5'h1c; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_79 = tableA_valid[29] ? _T_77 : 5'h1d; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_81 = tableA_valid[30] ? _T_79 : 5'h1e; // @[DFCTableA.scala 79:21]
  wire [4:0] _T_83 = tableA_valid[31] ? _T_81 : 5'h1f; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_85 = tableA_valid[32] ? {{1'd0}, _T_83} : 6'h20; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_87 = tableA_valid[33] ? _T_85 : 6'h21; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_89 = tableA_valid[34] ? _T_87 : 6'h22; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_91 = tableA_valid[35] ? _T_89 : 6'h23; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_93 = tableA_valid[36] ? _T_91 : 6'h24; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_95 = tableA_valid[37] ? _T_93 : 6'h25; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_97 = tableA_valid[38] ? _T_95 : 6'h26; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_99 = tableA_valid[39] ? _T_97 : 6'h27; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_101 = tableA_valid[40] ? _T_99 : 6'h28; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_103 = tableA_valid[41] ? _T_101 : 6'h29; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_105 = tableA_valid[42] ? _T_103 : 6'h2a; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_107 = tableA_valid[43] ? _T_105 : 6'h2b; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_109 = tableA_valid[44] ? _T_107 : 6'h2c; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_111 = tableA_valid[45] ? _T_109 : 6'h2d; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_113 = tableA_valid[46] ? _T_111 : 6'h2e; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_115 = tableA_valid[47] ? _T_113 : 6'h2f; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_117 = tableA_valid[48] ? _T_115 : 6'h30; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_119 = tableA_valid[49] ? _T_117 : 6'h31; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_121 = tableA_valid[50] ? _T_119 : 6'h32; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_123 = tableA_valid[51] ? _T_121 : 6'h33; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_125 = tableA_valid[52] ? _T_123 : 6'h34; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_127 = tableA_valid[53] ? _T_125 : 6'h35; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_129 = tableA_valid[54] ? _T_127 : 6'h36; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_131 = tableA_valid[55] ? _T_129 : 6'h37; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_133 = tableA_valid[56] ? _T_131 : 6'h38; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_135 = tableA_valid[57] ? _T_133 : 6'h39; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_137 = tableA_valid[58] ? _T_135 : 6'h3a; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_139 = tableA_valid[59] ? _T_137 : 6'h3b; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_141 = tableA_valid[60] ? _T_139 : 6'h3c; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_143 = tableA_valid[61] ? _T_141 : 6'h3d; // @[DFCTableA.scala 79:21]
  wire [5:0] _T_145 = tableA_valid[62] ? _T_143 : 6'h3e; // @[DFCTableA.scala 79:21]
  wire [5:0] empty_addr = tableA_valid[63] ? _T_145 : 6'h3f; // @[DFCTableA.scala 79:21]
  wire [1:0] _T_150 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_1_data ? 2'h2 : {{1'd0}, io_cpu_w_data_bits_wPid
     == infoMetaMem_pid_MPORT_data}; // @[DFCTableA.scala 84:21]
  wire [1:0] _T_152 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_2_data ? 2'h3 : _T_150; // @[DFCTableA.scala 84:21]
  wire [2:0] _T_154 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_3_data ? 3'h4 : {{1'd0}, _T_152}; // @[DFCTableA.scala 84:21]
  wire [2:0] _T_156 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_4_data ? 3'h5 : _T_154; // @[DFCTableA.scala 84:21]
  wire [2:0] _T_158 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_5_data ? 3'h6 : _T_156; // @[DFCTableA.scala 84:21]
  wire [2:0] _T_160 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_6_data ? 3'h7 : _T_158; // @[DFCTableA.scala 84:21]
  wire [3:0] _T_162 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_7_data ? 4'h8 : {{1'd0}, _T_160}; // @[DFCTableA.scala 84:21]
  wire [3:0] _T_164 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_8_data ? 4'h9 : _T_162; // @[DFCTableA.scala 84:21]
  wire [3:0] _T_166 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_9_data ? 4'ha : _T_164; // @[DFCTableA.scala 84:21]
  wire [3:0] _T_168 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_10_data ? 4'hb : _T_166; // @[DFCTableA.scala 84:21]
  wire [3:0] _T_170 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_11_data ? 4'hc : _T_168; // @[DFCTableA.scala 84:21]
  wire [3:0] _T_172 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_12_data ? 4'hd : _T_170; // @[DFCTableA.scala 84:21]
  wire [3:0] _T_174 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_13_data ? 4'he : _T_172; // @[DFCTableA.scala 84:21]
  wire [3:0] _T_176 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_14_data ? 4'hf : _T_174; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_178 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_15_data ? 5'h10 : {{1'd0}, _T_176}; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_180 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_16_data ? 5'h11 : _T_178; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_182 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_17_data ? 5'h12 : _T_180; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_184 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_18_data ? 5'h13 : _T_182; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_186 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_19_data ? 5'h14 : _T_184; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_188 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_20_data ? 5'h15 : _T_186; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_190 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_21_data ? 5'h16 : _T_188; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_192 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_22_data ? 5'h17 : _T_190; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_194 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_23_data ? 5'h18 : _T_192; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_196 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_24_data ? 5'h19 : _T_194; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_198 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_25_data ? 5'h1a : _T_196; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_200 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_26_data ? 5'h1b : _T_198; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_202 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_27_data ? 5'h1c : _T_200; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_204 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_28_data ? 5'h1d : _T_202; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_206 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_29_data ? 5'h1e : _T_204; // @[DFCTableA.scala 84:21]
  wire [4:0] _T_208 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_30_data ? 5'h1f : _T_206; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_210 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_31_data ? 6'h20 : {{1'd0}, _T_208}; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_212 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_32_data ? 6'h21 : _T_210; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_214 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_33_data ? 6'h22 : _T_212; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_216 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_34_data ? 6'h23 : _T_214; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_218 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_35_data ? 6'h24 : _T_216; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_220 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_36_data ? 6'h25 : _T_218; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_222 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_37_data ? 6'h26 : _T_220; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_224 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_38_data ? 6'h27 : _T_222; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_226 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_39_data ? 6'h28 : _T_224; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_228 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_40_data ? 6'h29 : _T_226; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_230 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_41_data ? 6'h2a : _T_228; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_232 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_42_data ? 6'h2b : _T_230; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_234 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_43_data ? 6'h2c : _T_232; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_236 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_44_data ? 6'h2d : _T_234; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_238 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_45_data ? 6'h2e : _T_236; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_240 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_46_data ? 6'h2f : _T_238; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_242 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_47_data ? 6'h30 : _T_240; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_244 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_48_data ? 6'h31 : _T_242; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_246 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_49_data ? 6'h32 : _T_244; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_248 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_50_data ? 6'h33 : _T_246; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_250 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_51_data ? 6'h34 : _T_248; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_252 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_52_data ? 6'h35 : _T_250; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_254 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_53_data ? 6'h36 : _T_252; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_256 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_54_data ? 6'h37 : _T_254; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_258 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_55_data ? 6'h38 : _T_256; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_260 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_56_data ? 6'h39 : _T_258; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_262 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_57_data ? 6'h3a : _T_260; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_264 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_58_data ? 6'h3b : _T_262; // @[DFCTableA.scala 84:21]
  wire [5:0] _T_266 = io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_59_data ? 6'h3c : _T_264; // @[DFCTableA.scala 84:21]
  reg [5:0] foundAddr; // @[Reg.scala 15:16]
  wire [63:0] _T_273 = tableA_valid >> foundAddr; // @[DFCTableA.scala 87:53]
  wire  notFound = foundAddr == 6'h0 | ~_T_273[0]; // @[DFCTableA.scala 87:37]
  wire  notEmpty = empty_addr == 6'h0 | empty_addr[5:3] == 3'h0; // @[DFCTableA.scala 88:38]
  wire  _T_281 = io_tableD_lresp_ready & io_tableD_lresp_valid; // @[Decoupled.scala 40:37]
  wire  _T_282 = state == 4'h2; // @[DFCTableA.scala 103:14]
  wire [7:0] _GEN_5 = 6'h0 == table_wId ? 8'h1 : counter_0; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_6 = 6'h1 == table_wId ? 8'h1 : counter_1; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_7 = 6'h2 == table_wId ? 8'h1 : counter_2; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_8 = 6'h3 == table_wId ? 8'h1 : counter_3; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_9 = 6'h4 == table_wId ? 8'h1 : counter_4; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_10 = 6'h5 == table_wId ? 8'h1 : counter_5; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_11 = 6'h6 == table_wId ? 8'h1 : counter_6; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_12 = 6'h7 == table_wId ? 8'h1 : counter_7; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_13 = 6'h8 == table_wId ? 8'h1 : counter_8; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_14 = 6'h9 == table_wId ? 8'h1 : counter_9; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_15 = 6'ha == table_wId ? 8'h1 : counter_10; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_16 = 6'hb == table_wId ? 8'h1 : counter_11; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_17 = 6'hc == table_wId ? 8'h1 : counter_12; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_18 = 6'hd == table_wId ? 8'h1 : counter_13; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_19 = 6'he == table_wId ? 8'h1 : counter_14; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_20 = 6'hf == table_wId ? 8'h1 : counter_15; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_21 = 6'h10 == table_wId ? 8'h1 : counter_16; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_22 = 6'h11 == table_wId ? 8'h1 : counter_17; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_23 = 6'h12 == table_wId ? 8'h1 : counter_18; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_24 = 6'h13 == table_wId ? 8'h1 : counter_19; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_25 = 6'h14 == table_wId ? 8'h1 : counter_20; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_26 = 6'h15 == table_wId ? 8'h1 : counter_21; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_27 = 6'h16 == table_wId ? 8'h1 : counter_22; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_28 = 6'h17 == table_wId ? 8'h1 : counter_23; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_29 = 6'h18 == table_wId ? 8'h1 : counter_24; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_30 = 6'h19 == table_wId ? 8'h1 : counter_25; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_31 = 6'h1a == table_wId ? 8'h1 : counter_26; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_32 = 6'h1b == table_wId ? 8'h1 : counter_27; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_33 = 6'h1c == table_wId ? 8'h1 : counter_28; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_34 = 6'h1d == table_wId ? 8'h1 : counter_29; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_35 = 6'h1e == table_wId ? 8'h1 : counter_30; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_36 = 6'h1f == table_wId ? 8'h1 : counter_31; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_37 = 6'h20 == table_wId ? 8'h1 : counter_32; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_38 = 6'h21 == table_wId ? 8'h1 : counter_33; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_39 = 6'h22 == table_wId ? 8'h1 : counter_34; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_40 = 6'h23 == table_wId ? 8'h1 : counter_35; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_41 = 6'h24 == table_wId ? 8'h1 : counter_36; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_42 = 6'h25 == table_wId ? 8'h1 : counter_37; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_43 = 6'h26 == table_wId ? 8'h1 : counter_38; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_44 = 6'h27 == table_wId ? 8'h1 : counter_39; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_45 = 6'h28 == table_wId ? 8'h1 : counter_40; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_46 = 6'h29 == table_wId ? 8'h1 : counter_41; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_47 = 6'h2a == table_wId ? 8'h1 : counter_42; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_48 = 6'h2b == table_wId ? 8'h1 : counter_43; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_49 = 6'h2c == table_wId ? 8'h1 : counter_44; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_50 = 6'h2d == table_wId ? 8'h1 : counter_45; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_51 = 6'h2e == table_wId ? 8'h1 : counter_46; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_52 = 6'h2f == table_wId ? 8'h1 : counter_47; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_53 = 6'h30 == table_wId ? 8'h1 : counter_48; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_54 = 6'h31 == table_wId ? 8'h1 : counter_49; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_55 = 6'h32 == table_wId ? 8'h1 : counter_50; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_56 = 6'h33 == table_wId ? 8'h1 : counter_51; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_57 = 6'h34 == table_wId ? 8'h1 : counter_52; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_58 = 6'h35 == table_wId ? 8'h1 : counter_53; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_59 = 6'h36 == table_wId ? 8'h1 : counter_54; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_60 = 6'h37 == table_wId ? 8'h1 : counter_55; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_61 = 6'h38 == table_wId ? 8'h1 : counter_56; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_62 = 6'h39 == table_wId ? 8'h1 : counter_57; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_63 = 6'h3a == table_wId ? 8'h1 : counter_58; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_64 = 6'h3b == table_wId ? 8'h1 : counter_59; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_65 = 6'h3c == table_wId ? 8'h1 : counter_60; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_66 = 6'h3d == table_wId ? 8'h1 : counter_61; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_67 = 6'h3e == table_wId ? 8'h1 : counter_62; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_68 = 6'h3f == table_wId ? 8'h1 : counter_63; // @[DFCTableA.scala 106:26 DFCTableA.scala 106:26 DFCTableA.scala 29:20]
  wire [63:0] _T_283 = 64'h1 << table_wId; // @[DFCTableA.scala 107:42]
  wire [63:0] _T_284 = tableA_valid | _T_283; // @[DFCTableA.scala 107:42]
  wire [63:0] _T_285 = ~tableA_valid; // @[DFCTableA.scala 107:42]
  wire [63:0] _T_286 = _T_285 | _T_283; // @[DFCTableA.scala 107:42]
  wire [63:0] _T_287 = ~_T_286; // @[DFCTableA.scala 107:42]
  wire  _T_290 = ~reset; // @[DFCTableA.scala 109:13]
  wire [7:0] _GEN_70 = 6'h1 == table_wId ? counter_1 : counter_0; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_71 = 6'h2 == table_wId ? counter_2 : _GEN_70; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_72 = 6'h3 == table_wId ? counter_3 : _GEN_71; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_73 = 6'h4 == table_wId ? counter_4 : _GEN_72; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_74 = 6'h5 == table_wId ? counter_5 : _GEN_73; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_75 = 6'h6 == table_wId ? counter_6 : _GEN_74; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_76 = 6'h7 == table_wId ? counter_7 : _GEN_75; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_77 = 6'h8 == table_wId ? counter_8 : _GEN_76; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_78 = 6'h9 == table_wId ? counter_9 : _GEN_77; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_79 = 6'ha == table_wId ? counter_10 : _GEN_78; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_80 = 6'hb == table_wId ? counter_11 : _GEN_79; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_81 = 6'hc == table_wId ? counter_12 : _GEN_80; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_82 = 6'hd == table_wId ? counter_13 : _GEN_81; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_83 = 6'he == table_wId ? counter_14 : _GEN_82; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_84 = 6'hf == table_wId ? counter_15 : _GEN_83; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_85 = 6'h10 == table_wId ? counter_16 : _GEN_84; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_86 = 6'h11 == table_wId ? counter_17 : _GEN_85; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_87 = 6'h12 == table_wId ? counter_18 : _GEN_86; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_88 = 6'h13 == table_wId ? counter_19 : _GEN_87; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_89 = 6'h14 == table_wId ? counter_20 : _GEN_88; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_90 = 6'h15 == table_wId ? counter_21 : _GEN_89; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_91 = 6'h16 == table_wId ? counter_22 : _GEN_90; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_92 = 6'h17 == table_wId ? counter_23 : _GEN_91; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_93 = 6'h18 == table_wId ? counter_24 : _GEN_92; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_94 = 6'h19 == table_wId ? counter_25 : _GEN_93; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_95 = 6'h1a == table_wId ? counter_26 : _GEN_94; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_96 = 6'h1b == table_wId ? counter_27 : _GEN_95; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_97 = 6'h1c == table_wId ? counter_28 : _GEN_96; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_98 = 6'h1d == table_wId ? counter_29 : _GEN_97; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_99 = 6'h1e == table_wId ? counter_30 : _GEN_98; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_100 = 6'h1f == table_wId ? counter_31 : _GEN_99; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_101 = 6'h20 == table_wId ? counter_32 : _GEN_100; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_102 = 6'h21 == table_wId ? counter_33 : _GEN_101; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_103 = 6'h22 == table_wId ? counter_34 : _GEN_102; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_104 = 6'h23 == table_wId ? counter_35 : _GEN_103; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_105 = 6'h24 == table_wId ? counter_36 : _GEN_104; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_106 = 6'h25 == table_wId ? counter_37 : _GEN_105; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_107 = 6'h26 == table_wId ? counter_38 : _GEN_106; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_108 = 6'h27 == table_wId ? counter_39 : _GEN_107; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_109 = 6'h28 == table_wId ? counter_40 : _GEN_108; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_110 = 6'h29 == table_wId ? counter_41 : _GEN_109; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_111 = 6'h2a == table_wId ? counter_42 : _GEN_110; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_112 = 6'h2b == table_wId ? counter_43 : _GEN_111; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_113 = 6'h2c == table_wId ? counter_44 : _GEN_112; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_114 = 6'h2d == table_wId ? counter_45 : _GEN_113; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_115 = 6'h2e == table_wId ? counter_46 : _GEN_114; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_116 = 6'h2f == table_wId ? counter_47 : _GEN_115; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_117 = 6'h30 == table_wId ? counter_48 : _GEN_116; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_118 = 6'h31 == table_wId ? counter_49 : _GEN_117; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_119 = 6'h32 == table_wId ? counter_50 : _GEN_118; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_120 = 6'h33 == table_wId ? counter_51 : _GEN_119; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_121 = 6'h34 == table_wId ? counter_52 : _GEN_120; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_122 = 6'h35 == table_wId ? counter_53 : _GEN_121; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_123 = 6'h36 == table_wId ? counter_54 : _GEN_122; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_124 = 6'h37 == table_wId ? counter_55 : _GEN_123; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_125 = 6'h38 == table_wId ? counter_56 : _GEN_124; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_126 = 6'h39 == table_wId ? counter_57 : _GEN_125; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_127 = 6'h3a == table_wId ? counter_58 : _GEN_126; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_128 = 6'h3b == table_wId ? counter_59 : _GEN_127; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_129 = 6'h3c == table_wId ? counter_60 : _GEN_128; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_130 = 6'h3d == table_wId ? counter_61 : _GEN_129; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_131 = 6'h3e == table_wId ? counter_62 : _GEN_130; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _GEN_132 = 6'h3f == table_wId ? counter_63 : _GEN_131; // @[DFCTableA.scala 112:48 DFCTableA.scala 112:48]
  wire [7:0] _T_294 = _GEN_132 + 8'h1; // @[DFCTableA.scala 112:48]
  wire [7:0] _GEN_133 = 6'h0 == table_wId ? _T_294 : counter_0; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_134 = 6'h1 == table_wId ? _T_294 : counter_1; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_135 = 6'h2 == table_wId ? _T_294 : counter_2; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_136 = 6'h3 == table_wId ? _T_294 : counter_3; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_137 = 6'h4 == table_wId ? _T_294 : counter_4; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_138 = 6'h5 == table_wId ? _T_294 : counter_5; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_139 = 6'h6 == table_wId ? _T_294 : counter_6; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_140 = 6'h7 == table_wId ? _T_294 : counter_7; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_141 = 6'h8 == table_wId ? _T_294 : counter_8; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_142 = 6'h9 == table_wId ? _T_294 : counter_9; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_143 = 6'ha == table_wId ? _T_294 : counter_10; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_144 = 6'hb == table_wId ? _T_294 : counter_11; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_145 = 6'hc == table_wId ? _T_294 : counter_12; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_146 = 6'hd == table_wId ? _T_294 : counter_13; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_147 = 6'he == table_wId ? _T_294 : counter_14; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_148 = 6'hf == table_wId ? _T_294 : counter_15; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_149 = 6'h10 == table_wId ? _T_294 : counter_16; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_150 = 6'h11 == table_wId ? _T_294 : counter_17; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_151 = 6'h12 == table_wId ? _T_294 : counter_18; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_152 = 6'h13 == table_wId ? _T_294 : counter_19; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_153 = 6'h14 == table_wId ? _T_294 : counter_20; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_154 = 6'h15 == table_wId ? _T_294 : counter_21; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_155 = 6'h16 == table_wId ? _T_294 : counter_22; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_156 = 6'h17 == table_wId ? _T_294 : counter_23; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_157 = 6'h18 == table_wId ? _T_294 : counter_24; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_158 = 6'h19 == table_wId ? _T_294 : counter_25; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_159 = 6'h1a == table_wId ? _T_294 : counter_26; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_160 = 6'h1b == table_wId ? _T_294 : counter_27; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_161 = 6'h1c == table_wId ? _T_294 : counter_28; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_162 = 6'h1d == table_wId ? _T_294 : counter_29; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_163 = 6'h1e == table_wId ? _T_294 : counter_30; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_164 = 6'h1f == table_wId ? _T_294 : counter_31; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_165 = 6'h20 == table_wId ? _T_294 : counter_32; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_166 = 6'h21 == table_wId ? _T_294 : counter_33; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_167 = 6'h22 == table_wId ? _T_294 : counter_34; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_168 = 6'h23 == table_wId ? _T_294 : counter_35; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_169 = 6'h24 == table_wId ? _T_294 : counter_36; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_170 = 6'h25 == table_wId ? _T_294 : counter_37; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_171 = 6'h26 == table_wId ? _T_294 : counter_38; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_172 = 6'h27 == table_wId ? _T_294 : counter_39; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_173 = 6'h28 == table_wId ? _T_294 : counter_40; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_174 = 6'h29 == table_wId ? _T_294 : counter_41; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_175 = 6'h2a == table_wId ? _T_294 : counter_42; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_176 = 6'h2b == table_wId ? _T_294 : counter_43; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_177 = 6'h2c == table_wId ? _T_294 : counter_44; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_178 = 6'h2d == table_wId ? _T_294 : counter_45; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_179 = 6'h2e == table_wId ? _T_294 : counter_46; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_180 = 6'h2f == table_wId ? _T_294 : counter_47; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_181 = 6'h30 == table_wId ? _T_294 : counter_48; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_182 = 6'h31 == table_wId ? _T_294 : counter_49; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_183 = 6'h32 == table_wId ? _T_294 : counter_50; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_184 = 6'h33 == table_wId ? _T_294 : counter_51; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_185 = 6'h34 == table_wId ? _T_294 : counter_52; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_186 = 6'h35 == table_wId ? _T_294 : counter_53; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_187 = 6'h36 == table_wId ? _T_294 : counter_54; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_188 = 6'h37 == table_wId ? _T_294 : counter_55; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_189 = 6'h38 == table_wId ? _T_294 : counter_56; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_190 = 6'h39 == table_wId ? _T_294 : counter_57; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_191 = 6'h3a == table_wId ? _T_294 : counter_58; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_192 = 6'h3b == table_wId ? _T_294 : counter_59; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_193 = 6'h3c == table_wId ? _T_294 : counter_60; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_194 = 6'h3d == table_wId ? _T_294 : counter_61; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_195 = 6'h3e == table_wId ? _T_294 : counter_62; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_196 = 6'h3f == table_wId ? _T_294 : counter_63; // @[DFCTableA.scala 112:26 DFCTableA.scala 112:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_202 = notFound ? _GEN_5 : _GEN_133; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_203 = notFound ? _GEN_6 : _GEN_134; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_204 = notFound ? _GEN_7 : _GEN_135; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_205 = notFound ? _GEN_8 : _GEN_136; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_206 = notFound ? _GEN_9 : _GEN_137; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_207 = notFound ? _GEN_10 : _GEN_138; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_208 = notFound ? _GEN_11 : _GEN_139; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_209 = notFound ? _GEN_12 : _GEN_140; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_210 = notFound ? _GEN_13 : _GEN_141; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_211 = notFound ? _GEN_14 : _GEN_142; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_212 = notFound ? _GEN_15 : _GEN_143; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_213 = notFound ? _GEN_16 : _GEN_144; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_214 = notFound ? _GEN_17 : _GEN_145; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_215 = notFound ? _GEN_18 : _GEN_146; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_216 = notFound ? _GEN_19 : _GEN_147; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_217 = notFound ? _GEN_20 : _GEN_148; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_218 = notFound ? _GEN_21 : _GEN_149; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_219 = notFound ? _GEN_22 : _GEN_150; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_220 = notFound ? _GEN_23 : _GEN_151; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_221 = notFound ? _GEN_24 : _GEN_152; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_222 = notFound ? _GEN_25 : _GEN_153; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_223 = notFound ? _GEN_26 : _GEN_154; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_224 = notFound ? _GEN_27 : _GEN_155; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_225 = notFound ? _GEN_28 : _GEN_156; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_226 = notFound ? _GEN_29 : _GEN_157; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_227 = notFound ? _GEN_30 : _GEN_158; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_228 = notFound ? _GEN_31 : _GEN_159; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_229 = notFound ? _GEN_32 : _GEN_160; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_230 = notFound ? _GEN_33 : _GEN_161; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_231 = notFound ? _GEN_34 : _GEN_162; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_232 = notFound ? _GEN_35 : _GEN_163; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_233 = notFound ? _GEN_36 : _GEN_164; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_234 = notFound ? _GEN_37 : _GEN_165; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_235 = notFound ? _GEN_38 : _GEN_166; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_236 = notFound ? _GEN_39 : _GEN_167; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_237 = notFound ? _GEN_40 : _GEN_168; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_238 = notFound ? _GEN_41 : _GEN_169; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_239 = notFound ? _GEN_42 : _GEN_170; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_240 = notFound ? _GEN_43 : _GEN_171; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_241 = notFound ? _GEN_44 : _GEN_172; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_242 = notFound ? _GEN_45 : _GEN_173; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_243 = notFound ? _GEN_46 : _GEN_174; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_244 = notFound ? _GEN_47 : _GEN_175; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_245 = notFound ? _GEN_48 : _GEN_176; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_246 = notFound ? _GEN_49 : _GEN_177; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_247 = notFound ? _GEN_50 : _GEN_178; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_248 = notFound ? _GEN_51 : _GEN_179; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_249 = notFound ? _GEN_52 : _GEN_180; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_250 = notFound ? _GEN_53 : _GEN_181; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_251 = notFound ? _GEN_54 : _GEN_182; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_252 = notFound ? _GEN_55 : _GEN_183; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_253 = notFound ? _GEN_56 : _GEN_184; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_254 = notFound ? _GEN_57 : _GEN_185; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_255 = notFound ? _GEN_58 : _GEN_186; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_256 = notFound ? _GEN_59 : _GEN_187; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_257 = notFound ? _GEN_60 : _GEN_188; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_258 = notFound ? _GEN_61 : _GEN_189; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_259 = notFound ? _GEN_62 : _GEN_190; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_260 = notFound ? _GEN_63 : _GEN_191; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_261 = notFound ? _GEN_64 : _GEN_192; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_262 = notFound ? _GEN_65 : _GEN_193; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_263 = notFound ? _GEN_66 : _GEN_194; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_264 = notFound ? _GEN_67 : _GEN_195; // @[DFCTableA.scala 104:19]
  wire [7:0] _GEN_265 = notFound ? _GEN_68 : _GEN_196; // @[DFCTableA.scala 104:19]
  wire  _GEN_269 = state == 4'h2 & notFound; // @[DFCTableA.scala 103:26 DFCTableA.scala 30:32]
  wire [7:0] _GEN_272 = state == 4'h2 ? _GEN_202 : counter_0; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_273 = state == 4'h2 ? _GEN_203 : counter_1; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_274 = state == 4'h2 ? _GEN_204 : counter_2; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_275 = state == 4'h2 ? _GEN_205 : counter_3; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_276 = state == 4'h2 ? _GEN_206 : counter_4; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_277 = state == 4'h2 ? _GEN_207 : counter_5; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_278 = state == 4'h2 ? _GEN_208 : counter_6; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_279 = state == 4'h2 ? _GEN_209 : counter_7; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_280 = state == 4'h2 ? _GEN_210 : counter_8; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_281 = state == 4'h2 ? _GEN_211 : counter_9; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_282 = state == 4'h2 ? _GEN_212 : counter_10; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_283 = state == 4'h2 ? _GEN_213 : counter_11; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_284 = state == 4'h2 ? _GEN_214 : counter_12; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_285 = state == 4'h2 ? _GEN_215 : counter_13; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_286 = state == 4'h2 ? _GEN_216 : counter_14; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_287 = state == 4'h2 ? _GEN_217 : counter_15; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_288 = state == 4'h2 ? _GEN_218 : counter_16; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_289 = state == 4'h2 ? _GEN_219 : counter_17; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_290 = state == 4'h2 ? _GEN_220 : counter_18; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_291 = state == 4'h2 ? _GEN_221 : counter_19; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_292 = state == 4'h2 ? _GEN_222 : counter_20; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_293 = state == 4'h2 ? _GEN_223 : counter_21; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_294 = state == 4'h2 ? _GEN_224 : counter_22; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_295 = state == 4'h2 ? _GEN_225 : counter_23; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_296 = state == 4'h2 ? _GEN_226 : counter_24; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_297 = state == 4'h2 ? _GEN_227 : counter_25; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_298 = state == 4'h2 ? _GEN_228 : counter_26; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_299 = state == 4'h2 ? _GEN_229 : counter_27; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_300 = state == 4'h2 ? _GEN_230 : counter_28; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_301 = state == 4'h2 ? _GEN_231 : counter_29; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_302 = state == 4'h2 ? _GEN_232 : counter_30; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_303 = state == 4'h2 ? _GEN_233 : counter_31; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_304 = state == 4'h2 ? _GEN_234 : counter_32; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_305 = state == 4'h2 ? _GEN_235 : counter_33; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_306 = state == 4'h2 ? _GEN_236 : counter_34; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_307 = state == 4'h2 ? _GEN_237 : counter_35; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_308 = state == 4'h2 ? _GEN_238 : counter_36; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_309 = state == 4'h2 ? _GEN_239 : counter_37; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_310 = state == 4'h2 ? _GEN_240 : counter_38; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_311 = state == 4'h2 ? _GEN_241 : counter_39; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_312 = state == 4'h2 ? _GEN_242 : counter_40; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_313 = state == 4'h2 ? _GEN_243 : counter_41; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_314 = state == 4'h2 ? _GEN_244 : counter_42; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_315 = state == 4'h2 ? _GEN_245 : counter_43; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_316 = state == 4'h2 ? _GEN_246 : counter_44; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_317 = state == 4'h2 ? _GEN_247 : counter_45; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_318 = state == 4'h2 ? _GEN_248 : counter_46; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_319 = state == 4'h2 ? _GEN_249 : counter_47; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_320 = state == 4'h2 ? _GEN_250 : counter_48; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_321 = state == 4'h2 ? _GEN_251 : counter_49; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_322 = state == 4'h2 ? _GEN_252 : counter_50; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_323 = state == 4'h2 ? _GEN_253 : counter_51; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_324 = state == 4'h2 ? _GEN_254 : counter_52; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_325 = state == 4'h2 ? _GEN_255 : counter_53; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_326 = state == 4'h2 ? _GEN_256 : counter_54; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_327 = state == 4'h2 ? _GEN_257 : counter_55; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_328 = state == 4'h2 ? _GEN_258 : counter_56; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_329 = state == 4'h2 ? _GEN_259 : counter_57; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_330 = state == 4'h2 ? _GEN_260 : counter_58; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_331 = state == 4'h2 ? _GEN_261 : counter_59; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_332 = state == 4'h2 ? _GEN_262 : counter_60; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_333 = state == 4'h2 ? _GEN_263 : counter_61; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_334 = state == 4'h2 ? _GEN_264 : counter_62; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire [7:0] _GEN_335 = state == 4'h2 ? _GEN_265 : counter_63; // @[DFCTableA.scala 103:26 DFCTableA.scala 29:20]
  wire  _T_301 = state == 4'h7 & _GEN_132 != 8'h1; // @[DFCTableA.scala 119:27]
  wire [7:0] _T_303 = _GEN_132 - 8'h1; // @[DFCTableA.scala 120:46]
  wire  _T_309 = state == 4'h8; // @[DFCTableA.scala 126:14]
  wire  _T_310 = laststate != 4'h8; // @[DFCTableA.scala 126:38]
  wire  _T_311 = state == 4'h8 & laststate != 4'h8; // @[DFCTableA.scala 126:25]
  wire  _T_323 = 4'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_324 = io_tableD_ldata_ready & io_tableD_ldata_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_476 = _T_324 ? 4'h6 : state; // @[DFCTableA.scala 144:37 DFCTableA.scala 145:17 DFCTableA.scala 34:22]
  wire [3:0] _GEN_478 = io_cpu_l_data_valid ? _GEN_476 : state; // @[DFCTableA.scala 142:38 DFCTableA.scala 34:22]
  wire  _GEN_480 = io_cpu_w_data_valid ? 1'h0 : io_cpu_l_data_valid; // @[DFCTableA.scala 140:32 DFCTableA.scala 59:25]
  wire  _T_325 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_326 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_327 = io_tableD_wdata_ready & io_tableD_wdata_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_481 = _T_327 ? 4'h3 : state; // @[DFCTableA.scala 154:35 DFCTableA.scala 155:15 DFCTableA.scala 34:22]
  wire  _T_328 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_329 = io_tableD_wresp_ready & io_tableD_wresp_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_482 = io_tableD_wresp_bits ? 4'h5 : 4'h0; // @[DFCTableA.scala 165:41 DFCTableA.scala 166:18 DFCTableA.scala 168:18]
  wire  _GEN_483 = notEmpty | full_a; // @[DFCTableA.scala 162:23 DFCTableA.scala 163:18 DFCTableA.scala 43:23]
  wire [3:0] _GEN_484 = notEmpty ? 4'h4 : _GEN_482; // @[DFCTableA.scala 162:23 DFCTableA.scala 164:18]
  wire  _GEN_485 = _T_329 ? io_tableD_wresp_bits : full_d; // @[DFCTableA.scala 160:35 DFCTableA.scala 161:16 DFCTableA.scala 45:23]
  wire  _GEN_486 = _T_329 ? _GEN_483 : full_a; // @[DFCTableA.scala 160:35 DFCTableA.scala 43:23]
  wire [3:0] _GEN_487 = _T_329 ? _GEN_484 : state; // @[DFCTableA.scala 160:35 DFCTableA.scala 34:22]
  wire  _T_330 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_488 = full_d ? 4'h5 : 4'h0; // @[DFCTableA.scala 179:29 DFCTableA.scala 180:19 DFCTableA.scala 182:19]
  wire [3:0] _GEN_489 = full_a ? 4'h4 : _GEN_488; // @[DFCTableA.scala 177:23 DFCTableA.scala 178:19]
  wire [3:0] _GEN_490 = io_tableD_lresp_bits_finish ? _GEN_489 : 4'h7; // @[DFCTableA.scala 176:42 DFCTableA.scala 185:17]
  wire [3:0] _GEN_491 = _T_281 ? _GEN_490 : state; // @[DFCTableA.scala 175:35 DFCTableA.scala 34:22]
  wire  _T_332 = 4'h7 == state; // @[Conditional.scala 37:30]
  wire  _GEN_492 = _GEN_132 == 8'h1 ? 1'h0 : full_a; // @[DFCTableA.scala 191:39 DFCTableA.scala 192:16 DFCTableA.scala 43:23]
  wire [3:0] _GEN_493 = _GEN_132 == 8'h1 ? 4'h8 : 4'h6; // @[DFCTableA.scala 191:39 DFCTableA.scala 193:15 DFCTableA.scala 195:15]
  wire  _T_334 = 4'h8 == state; // @[Conditional.scala 37:30]
  wire  _T_335 = io_cpu_expt_data_ready & io_cpu_expt_data_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_494 = _T_335 ? 4'h6 : state; // @[DFCTableA.scala 200:36 DFCTableA.scala 201:15 DFCTableA.scala 34:22]
  wire  _T_336 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_338 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_499 = _T_338 & io_cpu_l_data_valid; // @[Conditional.scala 39:67 DFCTableA.scala 59:25]
  wire [3:0] _GEN_500 = _T_338 ? _GEN_478 : state; // @[Conditional.scala 39:67 DFCTableA.scala 34:22]
  wire  _GEN_501 = _T_336 ? io_cpu_l_data_valid : _GEN_499; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_502 = _T_336 ? _GEN_478 : _GEN_500; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_504 = _T_334 ? _GEN_494 : _GEN_502; // @[Conditional.scala 39:67]
  wire  _GEN_505 = _T_334 ? 1'h0 : _GEN_501; // @[Conditional.scala 39:67 DFCTableA.scala 59:25]
  wire  _GEN_506 = _T_332 ? 1'h0 : full_d; // @[Conditional.scala 39:67 DFCTableA.scala 190:14 DFCTableA.scala 45:23]
  wire  _GEN_507 = _T_332 ? _GEN_492 : full_a; // @[Conditional.scala 39:67 DFCTableA.scala 43:23]
  wire [3:0] _GEN_508 = _T_332 ? _GEN_493 : _GEN_504; // @[Conditional.scala 39:67]
  wire  _GEN_509 = _T_332 ? 1'h0 : _T_334; // @[Conditional.scala 39:67 DFCTableA.scala 63:26]
  wire  _GEN_510 = _T_332 ? 1'h0 : _GEN_505; // @[Conditional.scala 39:67 DFCTableA.scala 59:25]
  wire [3:0] _GEN_512 = _T_330 ? _GEN_491 : _GEN_508; // @[Conditional.scala 39:67]
  wire  _GEN_513 = _T_330 ? full_d : _GEN_506; // @[Conditional.scala 39:67 DFCTableA.scala 45:23]
  wire  _GEN_514 = _T_330 ? full_a : _GEN_507; // @[Conditional.scala 39:67 DFCTableA.scala 43:23]
  wire  _GEN_515 = _T_330 ? 1'h0 : _GEN_509; // @[Conditional.scala 39:67 DFCTableA.scala 63:26]
  wire  _GEN_516 = _T_330 ? 1'h0 : _GEN_510; // @[Conditional.scala 39:67 DFCTableA.scala 59:25]
  wire  _GEN_518 = _T_328 ? _GEN_485 : _GEN_513; // @[Conditional.scala 39:67]
  wire  _GEN_519 = _T_328 ? _GEN_486 : _GEN_514; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_520 = _T_328 ? _GEN_487 : _GEN_512; // @[Conditional.scala 39:67]
  wire  _GEN_521 = _T_328 ? 1'h0 : _T_330; // @[Conditional.scala 39:67 DFCTableA.scala 61:25]
  wire  _GEN_522 = _T_328 ? 1'h0 : _GEN_515; // @[Conditional.scala 39:67 DFCTableA.scala 63:26]
  wire  _GEN_523 = _T_328 ? 1'h0 : _GEN_516; // @[Conditional.scala 39:67 DFCTableA.scala 59:25]
  wire  _GEN_526 = _T_326 ? 1'h0 : _T_328; // @[Conditional.scala 39:67 DFCTableA.scala 57:25]
  wire  _GEN_529 = _T_326 ? 1'h0 : _GEN_521; // @[Conditional.scala 39:67 DFCTableA.scala 61:25]
  wire  _GEN_530 = _T_326 ? 1'h0 : _GEN_522; // @[Conditional.scala 39:67 DFCTableA.scala 63:26]
  wire  _GEN_531 = _T_326 ? 1'h0 : _GEN_523; // @[Conditional.scala 39:67 DFCTableA.scala 59:25]
  wire  _GEN_533 = _T_325 ? 1'h0 : _T_326; // @[Conditional.scala 39:67 DFCTableA.scala 54:25]
  wire  _GEN_534 = _T_325 ? 1'h0 : _GEN_526; // @[Conditional.scala 39:67 DFCTableA.scala 57:25]
  wire  _GEN_537 = _T_325 ? 1'h0 : _GEN_529; // @[Conditional.scala 39:67 DFCTableA.scala 61:25]
  wire  _GEN_538 = _T_325 ? 1'h0 : _GEN_530; // @[Conditional.scala 39:67 DFCTableA.scala 63:26]
  wire  _GEN_539 = _T_325 ? 1'h0 : _GEN_531; // @[Conditional.scala 39:67 DFCTableA.scala 59:25]
  wire  _GEN_551 = _T_282 & ~notFound; // @[DFCTableA.scala 114:13]
  assign infoMetaMem_pid_MPORT_addr = 6'h1;
  assign infoMetaMem_pid_MPORT_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_1_addr = 6'h2;
  assign infoMetaMem_pid_MPORT_1_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_1_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_2_addr = 6'h3;
  assign infoMetaMem_pid_MPORT_2_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_2_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_3_addr = 6'h4;
  assign infoMetaMem_pid_MPORT_3_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_3_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_4_addr = 6'h5;
  assign infoMetaMem_pid_MPORT_4_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_4_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_5_addr = 6'h6;
  assign infoMetaMem_pid_MPORT_5_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_5_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_6_addr = 6'h7;
  assign infoMetaMem_pid_MPORT_6_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_6_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_7_addr = 6'h8;
  assign infoMetaMem_pid_MPORT_7_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_7_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_8_addr = 6'h9;
  assign infoMetaMem_pid_MPORT_8_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_8_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_9_addr = 6'ha;
  assign infoMetaMem_pid_MPORT_9_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_9_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_10_addr = 6'hb;
  assign infoMetaMem_pid_MPORT_10_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_10_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_11_addr = 6'hc;
  assign infoMetaMem_pid_MPORT_11_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_11_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_12_addr = 6'hd;
  assign infoMetaMem_pid_MPORT_12_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_12_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_13_addr = 6'he;
  assign infoMetaMem_pid_MPORT_13_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_13_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_14_addr = 6'hf;
  assign infoMetaMem_pid_MPORT_14_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_14_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_15_addr = 6'h10;
  assign infoMetaMem_pid_MPORT_15_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_15_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_16_addr = 6'h11;
  assign infoMetaMem_pid_MPORT_16_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_16_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_17_addr = 6'h12;
  assign infoMetaMem_pid_MPORT_17_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_17_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_18_addr = 6'h13;
  assign infoMetaMem_pid_MPORT_18_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_18_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_19_addr = 6'h14;
  assign infoMetaMem_pid_MPORT_19_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_19_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_20_addr = 6'h15;
  assign infoMetaMem_pid_MPORT_20_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_20_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_21_addr = 6'h16;
  assign infoMetaMem_pid_MPORT_21_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_21_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_22_addr = 6'h17;
  assign infoMetaMem_pid_MPORT_22_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_22_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_23_addr = 6'h18;
  assign infoMetaMem_pid_MPORT_23_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_23_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_24_addr = 6'h19;
  assign infoMetaMem_pid_MPORT_24_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_24_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_25_addr = 6'h1a;
  assign infoMetaMem_pid_MPORT_25_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_25_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_26_addr = 6'h1b;
  assign infoMetaMem_pid_MPORT_26_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_26_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_27_addr = 6'h1c;
  assign infoMetaMem_pid_MPORT_27_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_27_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_28_addr = 6'h1d;
  assign infoMetaMem_pid_MPORT_28_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_28_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_29_addr = 6'h1e;
  assign infoMetaMem_pid_MPORT_29_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_29_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_30_addr = 6'h1f;
  assign infoMetaMem_pid_MPORT_30_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_30_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_31_addr = 6'h20;
  assign infoMetaMem_pid_MPORT_31_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_31_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_32_addr = 6'h21;
  assign infoMetaMem_pid_MPORT_32_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_32_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_33_addr = 6'h22;
  assign infoMetaMem_pid_MPORT_33_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_33_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_34_addr = 6'h23;
  assign infoMetaMem_pid_MPORT_34_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_34_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_35_addr = 6'h24;
  assign infoMetaMem_pid_MPORT_35_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_35_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_36_addr = 6'h25;
  assign infoMetaMem_pid_MPORT_36_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_36_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_37_addr = 6'h26;
  assign infoMetaMem_pid_MPORT_37_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_37_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_38_addr = 6'h27;
  assign infoMetaMem_pid_MPORT_38_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_38_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_39_addr = 6'h28;
  assign infoMetaMem_pid_MPORT_39_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_39_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_40_addr = 6'h29;
  assign infoMetaMem_pid_MPORT_40_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_40_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_41_addr = 6'h2a;
  assign infoMetaMem_pid_MPORT_41_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_41_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_42_addr = 6'h2b;
  assign infoMetaMem_pid_MPORT_42_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_42_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_43_addr = 6'h2c;
  assign infoMetaMem_pid_MPORT_43_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_43_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_44_addr = 6'h2d;
  assign infoMetaMem_pid_MPORT_44_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_44_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_45_addr = 6'h2e;
  assign infoMetaMem_pid_MPORT_45_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_45_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_46_addr = 6'h2f;
  assign infoMetaMem_pid_MPORT_46_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_46_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_47_addr = 6'h30;
  assign infoMetaMem_pid_MPORT_47_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_47_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_48_addr = 6'h31;
  assign infoMetaMem_pid_MPORT_48_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_48_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_49_addr = 6'h32;
  assign infoMetaMem_pid_MPORT_49_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_49_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_50_addr = 6'h33;
  assign infoMetaMem_pid_MPORT_50_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_50_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_51_addr = 6'h34;
  assign infoMetaMem_pid_MPORT_51_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_51_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_52_addr = 6'h35;
  assign infoMetaMem_pid_MPORT_52_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_52_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_53_addr = 6'h36;
  assign infoMetaMem_pid_MPORT_53_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_53_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_54_addr = 6'h37;
  assign infoMetaMem_pid_MPORT_54_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_54_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_55_addr = 6'h38;
  assign infoMetaMem_pid_MPORT_55_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_55_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_56_addr = 6'h39;
  assign infoMetaMem_pid_MPORT_56_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_56_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_57_addr = 6'h3a;
  assign infoMetaMem_pid_MPORT_57_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_57_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_58_addr = 6'h3b;
  assign infoMetaMem_pid_MPORT_58_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_58_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_59_addr = 6'h3c;
  assign infoMetaMem_pid_MPORT_59_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_59_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_60_addr = 6'h3d;
  assign infoMetaMem_pid_MPORT_60_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_60_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_61_addr = 6'h3e;
  assign infoMetaMem_pid_MPORT_61_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_61_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_62_addr = 6'h3f;
  assign infoMetaMem_pid_MPORT_62_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_62_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_64_addr = infoMetaMem_pid_MPORT_64_addr_pipe_0;
  assign infoMetaMem_pid_MPORT_64_data = infoMetaMem_pid[infoMetaMem_pid_MPORT_64_addr]; // @[DFCTableA.scala 30:32]
  assign infoMetaMem_pid_MPORT_63_data = pid_reg;
  assign infoMetaMem_pid_MPORT_63_addr = table_wId;
  assign infoMetaMem_pid_MPORT_63_mask = 1'h1;
  assign infoMetaMem_pid_MPORT_63_en = _T_282 & notFound;
  assign infoMetaMem_pid_MPORT_65_data = 16'h0;
  assign infoMetaMem_pid_MPORT_65_addr = table_wId;
  assign infoMetaMem_pid_MPORT_65_mask = 1'h1;
  assign infoMetaMem_pid_MPORT_65_en = _T_309 & _T_310;
  assign io_cpu_w_data_ready = state == 4'h0; // @[DFCTableA.scala 36:23]
  assign io_cpu_l_data_ready = is_idle | state == 4'h4 | state == 4'h5; // @[DFCTableA.scala 52:56]
  assign io_tableD_wdata_valid = _T_323 ? 1'h0 : _GEN_533; // @[Conditional.scala 40:58 DFCTableA.scala 54:25]
  assign io_tableD_wdata_bits_listenAddr = laddr_reg; // @[DFCTableA.scala 55:35]
  assign io_tableD_wdata_bits_tableAId = table_wId; // @[DFCTableA.scala 56:33]
  assign io_tableD_ldata_valid = _T_323 ? _GEN_480 : _GEN_539; // @[Conditional.scala 40:58]
  assign io_tableD_ldata_bits_listenAddr = io_cpu_l_data_bits_listenAddr; // @[DFCTableA.scala 60:35]
  assign io_tableD_wresp_ready = _T_323 ? 1'h0 : _GEN_534; // @[Conditional.scala 40:58 DFCTableA.scala 57:25]
  assign io_tableD_lresp_ready = _T_323 ? 1'h0 : _GEN_537; // @[Conditional.scala 40:58 DFCTableA.scala 61:25]
  assign io_cpu_expt_data_valid = _T_323 ? 1'h0 : _GEN_538; // @[Conditional.scala 40:58 DFCTableA.scala 63:26]
  assign io_cpu_expt_data_bits_pid = laststate == 4'h8 ? pid_reg : pid_act; // @[DFCTableA.scala 64:35]
  assign io_dfc_full_data_valid = (full_a_last | full_d_last) & (~full_a & ~full_d) | _T_15; // @[DFCTableA.scala 66:84]
  assign io_dfc_full_data_bits_full_sig = _T_13 & _T_14; // @[DFCTableA.scala 68:68]
  always @(posedge clock) begin
    if(infoMetaMem_pid_MPORT_63_en & infoMetaMem_pid_MPORT_63_mask) begin
      infoMetaMem_pid[infoMetaMem_pid_MPORT_63_addr] <= infoMetaMem_pid_MPORT_63_data; // @[DFCTableA.scala 30:32]
    end
    if(infoMetaMem_pid_MPORT_65_en & infoMetaMem_pid_MPORT_65_mask) begin
      infoMetaMem_pid[infoMetaMem_pid_MPORT_65_addr] <= infoMetaMem_pid_MPORT_65_data; // @[DFCTableA.scala 30:32]
    end
    infoMetaMem_pid_MPORT_64_en_pipe_0 <= io_tableD_lresp_ready & io_tableD_lresp_valid;
    if (io_tableD_lresp_ready & io_tableD_lresp_valid) begin
      infoMetaMem_pid_MPORT_64_addr_pipe_0 <= io_tableD_lresp_bits_tableAId;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h0 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_0 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_0 <= _GEN_272;
      end
    end else begin
      counter_0 <= _GEN_272;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h1 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_1 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_1 <= _GEN_273;
      end
    end else begin
      counter_1 <= _GEN_273;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h2 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_2 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_2 <= _GEN_274;
      end
    end else begin
      counter_2 <= _GEN_274;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h3 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_3 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_3 <= _GEN_275;
      end
    end else begin
      counter_3 <= _GEN_275;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h4 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_4 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_4 <= _GEN_276;
      end
    end else begin
      counter_4 <= _GEN_276;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h5 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_5 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_5 <= _GEN_277;
      end
    end else begin
      counter_5 <= _GEN_277;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h6 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_6 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_6 <= _GEN_278;
      end
    end else begin
      counter_6 <= _GEN_278;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h7 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_7 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_7 <= _GEN_279;
      end
    end else begin
      counter_7 <= _GEN_279;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h8 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_8 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_8 <= _GEN_280;
      end
    end else begin
      counter_8 <= _GEN_280;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h9 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_9 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_9 <= _GEN_281;
      end
    end else begin
      counter_9 <= _GEN_281;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'ha == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_10 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_10 <= _GEN_282;
      end
    end else begin
      counter_10 <= _GEN_282;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'hb == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_11 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_11 <= _GEN_283;
      end
    end else begin
      counter_11 <= _GEN_283;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'hc == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_12 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_12 <= _GEN_284;
      end
    end else begin
      counter_12 <= _GEN_284;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'hd == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_13 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_13 <= _GEN_285;
      end
    end else begin
      counter_13 <= _GEN_285;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'he == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_14 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_14 <= _GEN_286;
      end
    end else begin
      counter_14 <= _GEN_286;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'hf == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_15 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_15 <= _GEN_287;
      end
    end else begin
      counter_15 <= _GEN_287;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h10 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_16 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_16 <= _GEN_288;
      end
    end else begin
      counter_16 <= _GEN_288;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h11 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_17 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_17 <= _GEN_289;
      end
    end else begin
      counter_17 <= _GEN_289;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h12 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_18 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_18 <= _GEN_290;
      end
    end else begin
      counter_18 <= _GEN_290;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h13 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_19 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_19 <= _GEN_291;
      end
    end else begin
      counter_19 <= _GEN_291;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h14 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_20 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_20 <= _GEN_292;
      end
    end else begin
      counter_20 <= _GEN_292;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h15 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_21 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_21 <= _GEN_293;
      end
    end else begin
      counter_21 <= _GEN_293;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h16 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_22 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_22 <= _GEN_294;
      end
    end else begin
      counter_22 <= _GEN_294;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h17 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_23 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_23 <= _GEN_295;
      end
    end else begin
      counter_23 <= _GEN_295;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h18 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_24 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_24 <= _GEN_296;
      end
    end else begin
      counter_24 <= _GEN_296;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h19 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_25 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_25 <= _GEN_297;
      end
    end else begin
      counter_25 <= _GEN_297;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h1a == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_26 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_26 <= _GEN_298;
      end
    end else begin
      counter_26 <= _GEN_298;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h1b == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_27 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_27 <= _GEN_299;
      end
    end else begin
      counter_27 <= _GEN_299;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h1c == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_28 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_28 <= _GEN_300;
      end
    end else begin
      counter_28 <= _GEN_300;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h1d == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_29 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_29 <= _GEN_301;
      end
    end else begin
      counter_29 <= _GEN_301;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h1e == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_30 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_30 <= _GEN_302;
      end
    end else begin
      counter_30 <= _GEN_302;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h1f == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_31 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_31 <= _GEN_303;
      end
    end else begin
      counter_31 <= _GEN_303;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h20 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_32 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_32 <= _GEN_304;
      end
    end else begin
      counter_32 <= _GEN_304;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h21 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_33 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_33 <= _GEN_305;
      end
    end else begin
      counter_33 <= _GEN_305;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h22 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_34 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_34 <= _GEN_306;
      end
    end else begin
      counter_34 <= _GEN_306;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h23 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_35 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_35 <= _GEN_307;
      end
    end else begin
      counter_35 <= _GEN_307;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h24 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_36 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_36 <= _GEN_308;
      end
    end else begin
      counter_36 <= _GEN_308;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h25 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_37 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_37 <= _GEN_309;
      end
    end else begin
      counter_37 <= _GEN_309;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h26 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_38 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_38 <= _GEN_310;
      end
    end else begin
      counter_38 <= _GEN_310;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h27 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_39 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_39 <= _GEN_311;
      end
    end else begin
      counter_39 <= _GEN_311;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h28 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_40 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_40 <= _GEN_312;
      end
    end else begin
      counter_40 <= _GEN_312;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h29 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_41 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_41 <= _GEN_313;
      end
    end else begin
      counter_41 <= _GEN_313;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h2a == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_42 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_42 <= _GEN_314;
      end
    end else begin
      counter_42 <= _GEN_314;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h2b == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_43 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_43 <= _GEN_315;
      end
    end else begin
      counter_43 <= _GEN_315;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h2c == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_44 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_44 <= _GEN_316;
      end
    end else begin
      counter_44 <= _GEN_316;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h2d == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_45 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_45 <= _GEN_317;
      end
    end else begin
      counter_45 <= _GEN_317;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h2e == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_46 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_46 <= _GEN_318;
      end
    end else begin
      counter_46 <= _GEN_318;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h2f == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_47 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_47 <= _GEN_319;
      end
    end else begin
      counter_47 <= _GEN_319;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h30 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_48 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_48 <= _GEN_320;
      end
    end else begin
      counter_48 <= _GEN_320;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h31 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_49 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_49 <= _GEN_321;
      end
    end else begin
      counter_49 <= _GEN_321;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h32 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_50 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_50 <= _GEN_322;
      end
    end else begin
      counter_50 <= _GEN_322;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h33 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_51 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_51 <= _GEN_323;
      end
    end else begin
      counter_51 <= _GEN_323;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h34 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_52 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_52 <= _GEN_324;
      end
    end else begin
      counter_52 <= _GEN_324;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h35 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_53 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_53 <= _GEN_325;
      end
    end else begin
      counter_53 <= _GEN_325;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h36 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_54 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_54 <= _GEN_326;
      end
    end else begin
      counter_54 <= _GEN_326;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h37 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_55 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_55 <= _GEN_327;
      end
    end else begin
      counter_55 <= _GEN_327;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h38 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_56 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_56 <= _GEN_328;
      end
    end else begin
      counter_56 <= _GEN_328;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h39 == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_57 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_57 <= _GEN_329;
      end
    end else begin
      counter_57 <= _GEN_329;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h3a == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_58 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_58 <= _GEN_330;
      end
    end else begin
      counter_58 <= _GEN_330;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h3b == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_59 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_59 <= _GEN_331;
      end
    end else begin
      counter_59 <= _GEN_331;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h3c == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_60 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_60 <= _GEN_332;
      end
    end else begin
      counter_60 <= _GEN_332;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h3d == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_61 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_61 <= _GEN_333;
      end
    end else begin
      counter_61 <= _GEN_333;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h3e == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_62 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_62 <= _GEN_334;
      end
    end else begin
      counter_62 <= _GEN_334;
    end
    if (state == 4'h7 & _GEN_132 != 8'h1) begin // @[DFCTableA.scala 119:57]
      if (6'h3f == table_wId) begin // @[DFCTableA.scala 120:24]
        counter_63 <= _T_303; // @[DFCTableA.scala 120:24]
      end else begin
        counter_63 <= _GEN_335;
      end
    end else begin
      counter_63 <= _GEN_335;
    end
    if (reset) begin // @[DFCTableA.scala 31:29]
      tableA_valid <= 64'h0; // @[DFCTableA.scala 31:29]
    end else if (_T_311) begin // @[DFCTableA.scala 130:49]
      tableA_valid <= _T_287; // @[DFCTableA.scala 132:18]
    end else if (state == 4'h2) begin // @[DFCTableA.scala 103:26]
      if (notFound) begin // @[DFCTableA.scala 104:19]
        tableA_valid <= _T_284; // @[DFCTableA.scala 107:20]
      end
    end
    if (reset) begin // @[DFCTableA.scala 34:22]
      state <= 4'h0; // @[DFCTableA.scala 34:22]
    end else if (_T_323) begin // @[Conditional.scala 40:58]
      if (io_cpu_w_data_valid) begin // @[DFCTableA.scala 140:32]
        state <= 4'h1; // @[DFCTableA.scala 141:15]
      end else if (io_cpu_l_data_valid) begin // @[DFCTableA.scala 142:38]
        state <= _GEN_476;
      end
    end else if (_T_325) begin // @[Conditional.scala 39:67]
      state <= 4'h2; // @[DFCTableA.scala 150:13]
    end else if (_T_326) begin // @[Conditional.scala 39:67]
      state <= _GEN_481;
    end else begin
      state <= _GEN_520;
    end
    laststate <= state; // @[DFCTableA.scala 35:26]
    if (reset) begin // @[DFCTableA.scala 39:26]
      laddr_reg <= 32'h0; // @[DFCTableA.scala 39:26]
    end else if (wEn) begin // @[DFCTableA.scala 71:12]
      laddr_reg <= io_cpu_w_data_bits_listenAddr; // @[DFCTableA.scala 72:15]
    end
    if (reset) begin // @[DFCTableA.scala 40:24]
      pid_reg <= 16'h0; // @[DFCTableA.scala 40:24]
    end else if (state == 4'h8 & laststate != 4'h8) begin // @[DFCTableA.scala 126:49]
      pid_reg <= pid_act; // @[DFCTableA.scala 127:13]
    end else if (wEn) begin // @[DFCTableA.scala 71:12]
      pid_reg <= io_cpu_w_data_bits_wPid; // @[DFCTableA.scala 73:13]
    end
    if (reset) begin // @[DFCTableA.scala 41:24]
      pid_act <= 16'h0; // @[DFCTableA.scala 41:24]
    end else begin
      pid_act <= infoMetaMem_pid_MPORT_64_data; // @[DFCTableA.scala 125:11]
    end
    if (reset) begin // @[DFCTableA.scala 42:26]
      table_wId <= 6'h1; // @[DFCTableA.scala 42:26]
    end else if (_T_281) begin // @[DFCTableA.scala 94:31]
      table_wId <= io_tableD_lresp_bits_tableAId; // @[DFCTableA.scala 95:15]
    end else if (state == 4'h1) begin // @[DFCTableA.scala 91:26]
      if (notFound) begin // @[DFCTableA.scala 92:21]
        table_wId <= empty_addr;
      end else begin
        table_wId <= foundAddr;
      end
    end
    if (reset) begin // @[DFCTableA.scala 43:23]
      full_a <= 1'h0; // @[DFCTableA.scala 43:23]
    end else if (!(_T_323)) begin // @[Conditional.scala 40:58]
      if (!(_T_325)) begin // @[Conditional.scala 39:67]
        if (!(_T_326)) begin // @[Conditional.scala 39:67]
          full_a <= _GEN_519;
        end
      end
    end
    full_a_last <= full_a; // @[DFCTableA.scala 44:28]
    if (reset) begin // @[DFCTableA.scala 45:23]
      full_d <= 1'h0; // @[DFCTableA.scala 45:23]
    end else if (!(_T_323)) begin // @[Conditional.scala 40:58]
      if (!(_T_325)) begin // @[Conditional.scala 39:67]
        if (!(_T_326)) begin // @[Conditional.scala 39:67]
          full_d <= _GEN_518;
        end
      end
    end
    full_d_last <= full_d; // @[DFCTableA.scala 46:28]
    if (wEn) begin // @[Reg.scala 16:19]
      if (io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_62_data) begin // @[DFCTableA.scala 84:21]
        foundAddr <= 6'h3f;
      end else if (io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_61_data) begin // @[DFCTableA.scala 84:21]
        foundAddr <= 6'h3e;
      end else if (io_cpu_w_data_bits_wPid == infoMetaMem_pid_MPORT_60_data) begin // @[DFCTableA.scala 84:21]
        foundAddr <= 6'h3d;
      end else begin
        foundAddr <= _T_266;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_269 & ~reset) begin
          $fwrite(32'h80000002,"[WTA](id: %d).infoMeta.pid = %d\n",table_wId,pid_reg); // @[DFCTableA.scala 109:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_269 & _T_290) begin
          $fwrite(32'h80000002,"[WC](id: %d).counter = %d\n",table_wId,1'h1); // @[DFCTableA.scala 110:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_282 & ~notFound & _T_290) begin
          $fwrite(32'h80000002,"[WTA_EXIST](id: %d).infoMeta.pid = %d\n",table_wId,pid_reg); // @[DFCTableA.scala 114:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_551 & _T_290) begin
          $fwrite(32'h80000002,"[WC](id: %d).counter = %d\n",table_wId,_GEN_132); // @[DFCTableA.scala 115:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_301 & _T_290) begin
          $fwrite(32'h80000002,"[WC_DOWN](id: %d).counter = %d\n",table_wId,_GEN_132); // @[DFCTableA.scala 121:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_311 & _T_290) begin
          $fwrite(32'h80000002,"[LTA](id: %d).infoMeta.pid Init!\n",table_wId); // @[DFCTableA.scala 134:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    infoMetaMem_pid[initvar] = _RAND_0[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  infoMetaMem_pid_MPORT_64_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  infoMetaMem_pid_MPORT_64_addr_pipe_0 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  counter_0 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  counter_1 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  counter_2 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  counter_3 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  counter_4 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  counter_5 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  counter_6 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  counter_7 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  counter_8 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  counter_9 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  counter_10 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  counter_11 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  counter_12 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  counter_13 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  counter_14 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  counter_15 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  counter_16 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  counter_17 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  counter_18 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  counter_19 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  counter_20 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  counter_21 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  counter_22 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  counter_23 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  counter_24 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  counter_25 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  counter_26 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  counter_27 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  counter_28 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  counter_29 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  counter_30 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  counter_31 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  counter_32 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  counter_33 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  counter_34 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  counter_35 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  counter_36 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  counter_37 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  counter_38 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  counter_39 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  counter_40 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  counter_41 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  counter_42 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  counter_43 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  counter_44 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  counter_45 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  counter_46 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  counter_47 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  counter_48 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  counter_49 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  counter_50 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  counter_51 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  counter_52 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  counter_53 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  counter_54 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  counter_55 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  counter_56 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  counter_57 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  counter_58 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  counter_59 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  counter_60 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  counter_61 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  counter_62 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  counter_63 = _RAND_66[7:0];
  _RAND_67 = {2{`RANDOM}};
  tableA_valid = _RAND_67[63:0];
  _RAND_68 = {1{`RANDOM}};
  state = _RAND_68[3:0];
  _RAND_69 = {1{`RANDOM}};
  laststate = _RAND_69[3:0];
  _RAND_70 = {1{`RANDOM}};
  laddr_reg = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  pid_reg = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  pid_act = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  table_wId = _RAND_73[5:0];
  _RAND_74 = {1{`RANDOM}};
  full_a = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  full_a_last = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  full_d = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  full_d_last = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  foundAddr = _RAND_78[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DFC_TableD(
  input         clock,
  input         reset,
  output        io_tableA_wdata_ready,
  input         io_tableA_wdata_valid,
  input  [31:0] io_tableA_wdata_bits_listenAddr,
  input  [5:0]  io_tableA_wdata_bits_tableAId,
  output        io_tableA_ldata_ready,
  input         io_tableA_ldata_valid,
  input  [31:0] io_tableA_ldata_bits_listenAddr,
  input         io_tableA_wresp_ready,
  output        io_tableA_wresp_valid,
  output        io_tableA_wresp_bits,
  input         io_tableA_lresp_ready,
  output        io_tableA_lresp_valid,
  output [5:0]  io_tableA_lresp_bits_tableAId,
  output        io_tableA_lresp_bits_finish
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [255:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] addrMetaMem_listenAddr [0:255]; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_1_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_1_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_2_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_2_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_3_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_3_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_4_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_4_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_5_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_5_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_6_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_6_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_7_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_7_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_8_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_8_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_9_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_9_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_10_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_10_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_11_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_11_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_12_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_12_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_13_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_13_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_14_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_14_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_15_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_15_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_16_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_16_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_17_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_17_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_18_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_18_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_19_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_19_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_20_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_20_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_21_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_21_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_22_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_22_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_23_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_23_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_24_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_24_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_25_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_25_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_26_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_26_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_27_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_27_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_28_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_28_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_29_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_29_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_30_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_30_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_31_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_31_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_32_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_32_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_33_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_33_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_34_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_34_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_35_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_35_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_36_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_36_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_37_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_37_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_38_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_38_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_39_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_39_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_40_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_40_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_41_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_41_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_42_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_42_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_43_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_43_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_44_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_44_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_45_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_45_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_46_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_46_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_47_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_47_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_48_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_48_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_49_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_49_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_50_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_50_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_51_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_51_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_52_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_52_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_53_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_53_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_54_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_54_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_55_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_55_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_56_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_56_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_57_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_57_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_58_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_58_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_59_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_59_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_60_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_60_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_61_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_61_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_62_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_62_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_63_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_63_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_64_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_64_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_65_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_65_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_66_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_66_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_67_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_67_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_68_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_68_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_69_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_69_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_70_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_70_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_71_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_71_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_72_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_72_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_73_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_73_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_74_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_74_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_75_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_75_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_76_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_76_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_77_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_77_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_78_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_78_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_79_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_79_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_80_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_80_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_81_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_81_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_82_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_82_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_83_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_83_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_84_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_84_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_85_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_85_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_86_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_86_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_87_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_87_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_88_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_88_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_89_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_89_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_90_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_90_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_91_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_91_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_92_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_92_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_93_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_93_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_94_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_94_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_95_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_95_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_96_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_96_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_97_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_97_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_98_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_98_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_99_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_99_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_100_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_100_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_101_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_101_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_102_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_102_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_103_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_103_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_104_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_104_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_105_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_105_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_106_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_106_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_107_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_107_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_108_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_108_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_109_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_109_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_110_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_110_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_111_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_111_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_112_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_112_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_113_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_113_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_114_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_114_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_115_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_115_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_116_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_116_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_117_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_117_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_118_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_118_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_119_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_119_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_120_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_120_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_121_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_121_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_122_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_122_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_123_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_123_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_124_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_124_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_125_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_125_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_126_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_126_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_127_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_127_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_128_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_128_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_129_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_129_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_130_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_130_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_131_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_131_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_132_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_132_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_133_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_133_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_134_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_134_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_135_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_135_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_136_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_136_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_137_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_137_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_138_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_138_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_139_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_139_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_140_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_140_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_141_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_141_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_142_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_142_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_143_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_143_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_144_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_144_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_145_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_145_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_146_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_146_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_147_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_147_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_148_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_148_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_149_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_149_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_150_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_150_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_151_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_151_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_152_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_152_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_153_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_153_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_154_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_154_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_155_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_155_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_156_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_156_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_157_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_157_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_158_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_158_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_159_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_159_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_160_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_160_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_161_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_161_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_162_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_162_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_163_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_163_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_164_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_164_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_165_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_165_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_166_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_166_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_167_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_167_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_168_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_168_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_169_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_169_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_170_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_170_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_171_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_171_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_172_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_172_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_173_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_173_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_174_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_174_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_175_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_175_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_176_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_176_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_177_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_177_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_178_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_178_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_179_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_179_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_180_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_180_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_181_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_181_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_182_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_182_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_183_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_183_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_184_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_184_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_185_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_185_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_186_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_186_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_187_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_187_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_188_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_188_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_189_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_189_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_190_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_190_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_191_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_191_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_192_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_192_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_193_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_193_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_194_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_194_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_195_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_195_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_196_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_196_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_197_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_197_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_198_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_198_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_199_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_199_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_200_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_200_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_201_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_201_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_202_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_202_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_203_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_203_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_204_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_204_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_205_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_205_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_206_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_206_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_207_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_207_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_208_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_208_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_209_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_209_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_210_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_210_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_211_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_211_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_212_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_212_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_213_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_213_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_214_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_214_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_215_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_215_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_216_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_216_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_217_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_217_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_218_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_218_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_219_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_219_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_220_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_220_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_221_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_221_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_222_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_222_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_223_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_223_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_224_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_224_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_225_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_225_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_226_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_226_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_227_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_227_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_228_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_228_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_229_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_229_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_230_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_230_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_231_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_231_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_232_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_232_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_233_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_233_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_234_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_234_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_235_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_235_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_236_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_236_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_237_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_237_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_238_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_238_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_239_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_239_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_240_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_240_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_241_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_241_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_242_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_242_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_243_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_243_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_244_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_244_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_245_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_245_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_246_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_246_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_247_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_247_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_248_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_248_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_249_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_249_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_250_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_250_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_251_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_251_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_252_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_252_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_253_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_253_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_254_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_254_addr; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_256_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_256_addr; // @[DFCTableD.scala 25:32]
  wire  addrMetaMem_listenAddr_MPORT_256_mask; // @[DFCTableD.scala 25:32]
  wire  addrMetaMem_listenAddr_MPORT_256_en; // @[DFCTableD.scala 25:32]
  wire [31:0] addrMetaMem_listenAddr_MPORT_258_data; // @[DFCTableD.scala 25:32]
  wire [7:0] addrMetaMem_listenAddr_MPORT_258_addr; // @[DFCTableD.scala 25:32]
  wire  addrMetaMem_listenAddr_MPORT_258_mask; // @[DFCTableD.scala 25:32]
  wire  addrMetaMem_listenAddr_MPORT_258_en; // @[DFCTableD.scala 25:32]
  reg [5:0] infoMetaMem_tableAid [0:255]; // @[DFCTableD.scala 26:32]
  wire [5:0] infoMetaMem_tableAid_MPORT_255_data; // @[DFCTableD.scala 26:32]
  wire [7:0] infoMetaMem_tableAid_MPORT_255_addr; // @[DFCTableD.scala 26:32]
  wire [5:0] infoMetaMem_tableAid_MPORT_257_data; // @[DFCTableD.scala 26:32]
  wire [7:0] infoMetaMem_tableAid_MPORT_257_addr; // @[DFCTableD.scala 26:32]
  wire  infoMetaMem_tableAid_MPORT_257_mask; // @[DFCTableD.scala 26:32]
  wire  infoMetaMem_tableAid_MPORT_257_en; // @[DFCTableD.scala 26:32]
  wire [5:0] infoMetaMem_tableAid_MPORT_259_data; // @[DFCTableD.scala 26:32]
  wire [7:0] infoMetaMem_tableAid_MPORT_259_addr; // @[DFCTableD.scala 26:32]
  wire  infoMetaMem_tableAid_MPORT_259_mask; // @[DFCTableD.scala 26:32]
  wire  infoMetaMem_tableAid_MPORT_259_en; // @[DFCTableD.scala 26:32]
  reg [7:0] infoMetaMem_tableAid_MPORT_255_addr_pipe_0;
  reg [255:0] tableD_valid; // @[DFCTableD.scala 27:29]
  reg [2:0] state; // @[DFCTableD.scala 30:22]
  reg [2:0] laststate; // @[DFCTableD.scala 31:26]
  wire  is_idle = state == 3'h0; // @[DFCTableD.scala 32:23]
  reg [31:0] laddr_reg; // @[DFCTableD.scala 35:26]
  reg [5:0] tableAid_reg; // @[DFCTableD.scala 36:29]
  reg [7:0] tableD_Id; // @[DFCTableD.scala 37:26]
  reg [7:0] match_Id; // @[DFCTableD.scala 38:25]
  reg [5:0] cDown_Id; // @[DFCTableD.scala 39:25]
  reg [5:0] cDown_Id_reg; // @[DFCTableD.scala 40:29]
  wire  _T = state == 3'h5; // @[DFCTableD.scala 41:28]
  wire  _T_7 = tableD_valid[1] ? 1'h0 : 1'h1; // @[DFCTableD.scala 57:21]
  wire [1:0] _T_9 = tableD_valid[2] ? {{1'd0}, _T_7} : 2'h2; // @[DFCTableD.scala 57:21]
  wire [1:0] _T_11 = tableD_valid[3] ? _T_9 : 2'h3; // @[DFCTableD.scala 57:21]
  wire [2:0] _T_13 = tableD_valid[4] ? {{1'd0}, _T_11} : 3'h4; // @[DFCTableD.scala 57:21]
  wire [2:0] _T_15 = tableD_valid[5] ? _T_13 : 3'h5; // @[DFCTableD.scala 57:21]
  wire [2:0] _T_17 = tableD_valid[6] ? _T_15 : 3'h6; // @[DFCTableD.scala 57:21]
  wire [2:0] _T_19 = tableD_valid[7] ? _T_17 : 3'h7; // @[DFCTableD.scala 57:21]
  wire [3:0] _T_21 = tableD_valid[8] ? {{1'd0}, _T_19} : 4'h8; // @[DFCTableD.scala 57:21]
  wire [3:0] _T_23 = tableD_valid[9] ? _T_21 : 4'h9; // @[DFCTableD.scala 57:21]
  wire [3:0] _T_25 = tableD_valid[10] ? _T_23 : 4'ha; // @[DFCTableD.scala 57:21]
  wire [3:0] _T_27 = tableD_valid[11] ? _T_25 : 4'hb; // @[DFCTableD.scala 57:21]
  wire [3:0] _T_29 = tableD_valid[12] ? _T_27 : 4'hc; // @[DFCTableD.scala 57:21]
  wire [3:0] _T_31 = tableD_valid[13] ? _T_29 : 4'hd; // @[DFCTableD.scala 57:21]
  wire [3:0] _T_33 = tableD_valid[14] ? _T_31 : 4'he; // @[DFCTableD.scala 57:21]
  wire [3:0] _T_35 = tableD_valid[15] ? _T_33 : 4'hf; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_37 = tableD_valid[16] ? {{1'd0}, _T_35} : 5'h10; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_39 = tableD_valid[17] ? _T_37 : 5'h11; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_41 = tableD_valid[18] ? _T_39 : 5'h12; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_43 = tableD_valid[19] ? _T_41 : 5'h13; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_45 = tableD_valid[20] ? _T_43 : 5'h14; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_47 = tableD_valid[21] ? _T_45 : 5'h15; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_49 = tableD_valid[22] ? _T_47 : 5'h16; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_51 = tableD_valid[23] ? _T_49 : 5'h17; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_53 = tableD_valid[24] ? _T_51 : 5'h18; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_55 = tableD_valid[25] ? _T_53 : 5'h19; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_57 = tableD_valid[26] ? _T_55 : 5'h1a; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_59 = tableD_valid[27] ? _T_57 : 5'h1b; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_61 = tableD_valid[28] ? _T_59 : 5'h1c; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_63 = tableD_valid[29] ? _T_61 : 5'h1d; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_65 = tableD_valid[30] ? _T_63 : 5'h1e; // @[DFCTableD.scala 57:21]
  wire [4:0] _T_67 = tableD_valid[31] ? _T_65 : 5'h1f; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_69 = tableD_valid[32] ? {{1'd0}, _T_67} : 6'h20; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_71 = tableD_valid[33] ? _T_69 : 6'h21; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_73 = tableD_valid[34] ? _T_71 : 6'h22; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_75 = tableD_valid[35] ? _T_73 : 6'h23; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_77 = tableD_valid[36] ? _T_75 : 6'h24; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_79 = tableD_valid[37] ? _T_77 : 6'h25; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_81 = tableD_valid[38] ? _T_79 : 6'h26; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_83 = tableD_valid[39] ? _T_81 : 6'h27; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_85 = tableD_valid[40] ? _T_83 : 6'h28; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_87 = tableD_valid[41] ? _T_85 : 6'h29; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_89 = tableD_valid[42] ? _T_87 : 6'h2a; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_91 = tableD_valid[43] ? _T_89 : 6'h2b; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_93 = tableD_valid[44] ? _T_91 : 6'h2c; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_95 = tableD_valid[45] ? _T_93 : 6'h2d; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_97 = tableD_valid[46] ? _T_95 : 6'h2e; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_99 = tableD_valid[47] ? _T_97 : 6'h2f; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_101 = tableD_valid[48] ? _T_99 : 6'h30; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_103 = tableD_valid[49] ? _T_101 : 6'h31; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_105 = tableD_valid[50] ? _T_103 : 6'h32; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_107 = tableD_valid[51] ? _T_105 : 6'h33; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_109 = tableD_valid[52] ? _T_107 : 6'h34; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_111 = tableD_valid[53] ? _T_109 : 6'h35; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_113 = tableD_valid[54] ? _T_111 : 6'h36; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_115 = tableD_valid[55] ? _T_113 : 6'h37; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_117 = tableD_valid[56] ? _T_115 : 6'h38; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_119 = tableD_valid[57] ? _T_117 : 6'h39; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_121 = tableD_valid[58] ? _T_119 : 6'h3a; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_123 = tableD_valid[59] ? _T_121 : 6'h3b; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_125 = tableD_valid[60] ? _T_123 : 6'h3c; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_127 = tableD_valid[61] ? _T_125 : 6'h3d; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_129 = tableD_valid[62] ? _T_127 : 6'h3e; // @[DFCTableD.scala 57:21]
  wire [5:0] _T_131 = tableD_valid[63] ? _T_129 : 6'h3f; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_133 = tableD_valid[64] ? {{1'd0}, _T_131} : 7'h40; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_135 = tableD_valid[65] ? _T_133 : 7'h41; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_137 = tableD_valid[66] ? _T_135 : 7'h42; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_139 = tableD_valid[67] ? _T_137 : 7'h43; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_141 = tableD_valid[68] ? _T_139 : 7'h44; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_143 = tableD_valid[69] ? _T_141 : 7'h45; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_145 = tableD_valid[70] ? _T_143 : 7'h46; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_147 = tableD_valid[71] ? _T_145 : 7'h47; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_149 = tableD_valid[72] ? _T_147 : 7'h48; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_151 = tableD_valid[73] ? _T_149 : 7'h49; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_153 = tableD_valid[74] ? _T_151 : 7'h4a; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_155 = tableD_valid[75] ? _T_153 : 7'h4b; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_157 = tableD_valid[76] ? _T_155 : 7'h4c; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_159 = tableD_valid[77] ? _T_157 : 7'h4d; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_161 = tableD_valid[78] ? _T_159 : 7'h4e; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_163 = tableD_valid[79] ? _T_161 : 7'h4f; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_165 = tableD_valid[80] ? _T_163 : 7'h50; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_167 = tableD_valid[81] ? _T_165 : 7'h51; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_169 = tableD_valid[82] ? _T_167 : 7'h52; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_171 = tableD_valid[83] ? _T_169 : 7'h53; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_173 = tableD_valid[84] ? _T_171 : 7'h54; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_175 = tableD_valid[85] ? _T_173 : 7'h55; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_177 = tableD_valid[86] ? _T_175 : 7'h56; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_179 = tableD_valid[87] ? _T_177 : 7'h57; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_181 = tableD_valid[88] ? _T_179 : 7'h58; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_183 = tableD_valid[89] ? _T_181 : 7'h59; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_185 = tableD_valid[90] ? _T_183 : 7'h5a; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_187 = tableD_valid[91] ? _T_185 : 7'h5b; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_189 = tableD_valid[92] ? _T_187 : 7'h5c; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_191 = tableD_valid[93] ? _T_189 : 7'h5d; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_193 = tableD_valid[94] ? _T_191 : 7'h5e; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_195 = tableD_valid[95] ? _T_193 : 7'h5f; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_197 = tableD_valid[96] ? _T_195 : 7'h60; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_199 = tableD_valid[97] ? _T_197 : 7'h61; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_201 = tableD_valid[98] ? _T_199 : 7'h62; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_203 = tableD_valid[99] ? _T_201 : 7'h63; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_205 = tableD_valid[100] ? _T_203 : 7'h64; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_207 = tableD_valid[101] ? _T_205 : 7'h65; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_209 = tableD_valid[102] ? _T_207 : 7'h66; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_211 = tableD_valid[103] ? _T_209 : 7'h67; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_213 = tableD_valid[104] ? _T_211 : 7'h68; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_215 = tableD_valid[105] ? _T_213 : 7'h69; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_217 = tableD_valid[106] ? _T_215 : 7'h6a; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_219 = tableD_valid[107] ? _T_217 : 7'h6b; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_221 = tableD_valid[108] ? _T_219 : 7'h6c; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_223 = tableD_valid[109] ? _T_221 : 7'h6d; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_225 = tableD_valid[110] ? _T_223 : 7'h6e; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_227 = tableD_valid[111] ? _T_225 : 7'h6f; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_229 = tableD_valid[112] ? _T_227 : 7'h70; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_231 = tableD_valid[113] ? _T_229 : 7'h71; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_233 = tableD_valid[114] ? _T_231 : 7'h72; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_235 = tableD_valid[115] ? _T_233 : 7'h73; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_237 = tableD_valid[116] ? _T_235 : 7'h74; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_239 = tableD_valid[117] ? _T_237 : 7'h75; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_241 = tableD_valid[118] ? _T_239 : 7'h76; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_243 = tableD_valid[119] ? _T_241 : 7'h77; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_245 = tableD_valid[120] ? _T_243 : 7'h78; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_247 = tableD_valid[121] ? _T_245 : 7'h79; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_249 = tableD_valid[122] ? _T_247 : 7'h7a; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_251 = tableD_valid[123] ? _T_249 : 7'h7b; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_253 = tableD_valid[124] ? _T_251 : 7'h7c; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_255 = tableD_valid[125] ? _T_253 : 7'h7d; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_257 = tableD_valid[126] ? _T_255 : 7'h7e; // @[DFCTableD.scala 57:21]
  wire [6:0] _T_259 = tableD_valid[127] ? _T_257 : 7'h7f; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_261 = tableD_valid[128] ? {{1'd0}, _T_259} : 8'h80; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_263 = tableD_valid[129] ? _T_261 : 8'h81; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_265 = tableD_valid[130] ? _T_263 : 8'h82; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_267 = tableD_valid[131] ? _T_265 : 8'h83; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_269 = tableD_valid[132] ? _T_267 : 8'h84; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_271 = tableD_valid[133] ? _T_269 : 8'h85; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_273 = tableD_valid[134] ? _T_271 : 8'h86; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_275 = tableD_valid[135] ? _T_273 : 8'h87; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_277 = tableD_valid[136] ? _T_275 : 8'h88; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_279 = tableD_valid[137] ? _T_277 : 8'h89; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_281 = tableD_valid[138] ? _T_279 : 8'h8a; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_283 = tableD_valid[139] ? _T_281 : 8'h8b; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_285 = tableD_valid[140] ? _T_283 : 8'h8c; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_287 = tableD_valid[141] ? _T_285 : 8'h8d; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_289 = tableD_valid[142] ? _T_287 : 8'h8e; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_291 = tableD_valid[143] ? _T_289 : 8'h8f; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_293 = tableD_valid[144] ? _T_291 : 8'h90; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_295 = tableD_valid[145] ? _T_293 : 8'h91; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_297 = tableD_valid[146] ? _T_295 : 8'h92; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_299 = tableD_valid[147] ? _T_297 : 8'h93; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_301 = tableD_valid[148] ? _T_299 : 8'h94; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_303 = tableD_valid[149] ? _T_301 : 8'h95; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_305 = tableD_valid[150] ? _T_303 : 8'h96; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_307 = tableD_valid[151] ? _T_305 : 8'h97; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_309 = tableD_valid[152] ? _T_307 : 8'h98; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_311 = tableD_valid[153] ? _T_309 : 8'h99; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_313 = tableD_valid[154] ? _T_311 : 8'h9a; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_315 = tableD_valid[155] ? _T_313 : 8'h9b; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_317 = tableD_valid[156] ? _T_315 : 8'h9c; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_319 = tableD_valid[157] ? _T_317 : 8'h9d; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_321 = tableD_valid[158] ? _T_319 : 8'h9e; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_323 = tableD_valid[159] ? _T_321 : 8'h9f; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_325 = tableD_valid[160] ? _T_323 : 8'ha0; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_327 = tableD_valid[161] ? _T_325 : 8'ha1; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_329 = tableD_valid[162] ? _T_327 : 8'ha2; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_331 = tableD_valid[163] ? _T_329 : 8'ha3; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_333 = tableD_valid[164] ? _T_331 : 8'ha4; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_335 = tableD_valid[165] ? _T_333 : 8'ha5; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_337 = tableD_valid[166] ? _T_335 : 8'ha6; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_339 = tableD_valid[167] ? _T_337 : 8'ha7; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_341 = tableD_valid[168] ? _T_339 : 8'ha8; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_343 = tableD_valid[169] ? _T_341 : 8'ha9; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_345 = tableD_valid[170] ? _T_343 : 8'haa; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_347 = tableD_valid[171] ? _T_345 : 8'hab; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_349 = tableD_valid[172] ? _T_347 : 8'hac; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_351 = tableD_valid[173] ? _T_349 : 8'had; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_353 = tableD_valid[174] ? _T_351 : 8'hae; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_355 = tableD_valid[175] ? _T_353 : 8'haf; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_357 = tableD_valid[176] ? _T_355 : 8'hb0; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_359 = tableD_valid[177] ? _T_357 : 8'hb1; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_361 = tableD_valid[178] ? _T_359 : 8'hb2; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_363 = tableD_valid[179] ? _T_361 : 8'hb3; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_365 = tableD_valid[180] ? _T_363 : 8'hb4; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_367 = tableD_valid[181] ? _T_365 : 8'hb5; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_369 = tableD_valid[182] ? _T_367 : 8'hb6; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_371 = tableD_valid[183] ? _T_369 : 8'hb7; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_373 = tableD_valid[184] ? _T_371 : 8'hb8; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_375 = tableD_valid[185] ? _T_373 : 8'hb9; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_377 = tableD_valid[186] ? _T_375 : 8'hba; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_379 = tableD_valid[187] ? _T_377 : 8'hbb; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_381 = tableD_valid[188] ? _T_379 : 8'hbc; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_383 = tableD_valid[189] ? _T_381 : 8'hbd; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_385 = tableD_valid[190] ? _T_383 : 8'hbe; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_387 = tableD_valid[191] ? _T_385 : 8'hbf; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_389 = tableD_valid[192] ? _T_387 : 8'hc0; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_391 = tableD_valid[193] ? _T_389 : 8'hc1; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_393 = tableD_valid[194] ? _T_391 : 8'hc2; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_395 = tableD_valid[195] ? _T_393 : 8'hc3; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_397 = tableD_valid[196] ? _T_395 : 8'hc4; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_399 = tableD_valid[197] ? _T_397 : 8'hc5; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_401 = tableD_valid[198] ? _T_399 : 8'hc6; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_403 = tableD_valid[199] ? _T_401 : 8'hc7; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_405 = tableD_valid[200] ? _T_403 : 8'hc8; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_407 = tableD_valid[201] ? _T_405 : 8'hc9; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_409 = tableD_valid[202] ? _T_407 : 8'hca; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_411 = tableD_valid[203] ? _T_409 : 8'hcb; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_413 = tableD_valid[204] ? _T_411 : 8'hcc; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_415 = tableD_valid[205] ? _T_413 : 8'hcd; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_417 = tableD_valid[206] ? _T_415 : 8'hce; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_419 = tableD_valid[207] ? _T_417 : 8'hcf; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_421 = tableD_valid[208] ? _T_419 : 8'hd0; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_423 = tableD_valid[209] ? _T_421 : 8'hd1; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_425 = tableD_valid[210] ? _T_423 : 8'hd2; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_427 = tableD_valid[211] ? _T_425 : 8'hd3; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_429 = tableD_valid[212] ? _T_427 : 8'hd4; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_431 = tableD_valid[213] ? _T_429 : 8'hd5; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_433 = tableD_valid[214] ? _T_431 : 8'hd6; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_435 = tableD_valid[215] ? _T_433 : 8'hd7; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_437 = tableD_valid[216] ? _T_435 : 8'hd8; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_439 = tableD_valid[217] ? _T_437 : 8'hd9; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_441 = tableD_valid[218] ? _T_439 : 8'hda; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_443 = tableD_valid[219] ? _T_441 : 8'hdb; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_445 = tableD_valid[220] ? _T_443 : 8'hdc; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_447 = tableD_valid[221] ? _T_445 : 8'hdd; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_449 = tableD_valid[222] ? _T_447 : 8'hde; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_451 = tableD_valid[223] ? _T_449 : 8'hdf; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_453 = tableD_valid[224] ? _T_451 : 8'he0; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_455 = tableD_valid[225] ? _T_453 : 8'he1; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_457 = tableD_valid[226] ? _T_455 : 8'he2; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_459 = tableD_valid[227] ? _T_457 : 8'he3; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_461 = tableD_valid[228] ? _T_459 : 8'he4; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_463 = tableD_valid[229] ? _T_461 : 8'he5; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_465 = tableD_valid[230] ? _T_463 : 8'he6; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_467 = tableD_valid[231] ? _T_465 : 8'he7; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_469 = tableD_valid[232] ? _T_467 : 8'he8; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_471 = tableD_valid[233] ? _T_469 : 8'he9; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_473 = tableD_valid[234] ? _T_471 : 8'hea; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_475 = tableD_valid[235] ? _T_473 : 8'heb; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_477 = tableD_valid[236] ? _T_475 : 8'hec; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_479 = tableD_valid[237] ? _T_477 : 8'hed; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_481 = tableD_valid[238] ? _T_479 : 8'hee; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_483 = tableD_valid[239] ? _T_481 : 8'hef; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_485 = tableD_valid[240] ? _T_483 : 8'hf0; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_487 = tableD_valid[241] ? _T_485 : 8'hf1; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_489 = tableD_valid[242] ? _T_487 : 8'hf2; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_491 = tableD_valid[243] ? _T_489 : 8'hf3; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_493 = tableD_valid[244] ? _T_491 : 8'hf4; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_495 = tableD_valid[245] ? _T_493 : 8'hf5; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_497 = tableD_valid[246] ? _T_495 : 8'hf6; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_499 = tableD_valid[247] ? _T_497 : 8'hf7; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_501 = tableD_valid[248] ? _T_499 : 8'hf8; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_503 = tableD_valid[249] ? _T_501 : 8'hf9; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_505 = tableD_valid[250] ? _T_503 : 8'hfa; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_507 = tableD_valid[251] ? _T_505 : 8'hfb; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_509 = tableD_valid[252] ? _T_507 : 8'hfc; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_511 = tableD_valid[253] ? _T_509 : 8'hfd; // @[DFCTableD.scala 57:21]
  wire [7:0] _T_513 = tableD_valid[254] ? _T_511 : 8'hfe; // @[DFCTableD.scala 57:21]
  wire [7:0] empty_addr = tableD_valid[255] ? _T_513 : 8'hff; // @[DFCTableD.scala 57:21]
  wire  notEmpty = empty_addr == 8'h0 | empty_addr[7:3] == 5'h0; // @[DFCTableD.scala 59:38]
  wire [1:0] _T_523 = laddr_reg == addrMetaMem_listenAddr_MPORT_1_data ? 2'h2 : {{1'd0}, laddr_reg ==
    addrMetaMem_listenAddr_MPORT_data}; // @[DFCTableD.scala 72:21]
  wire [1:0] _T_525 = laddr_reg == addrMetaMem_listenAddr_MPORT_2_data ? 2'h3 : _T_523; // @[DFCTableD.scala 72:21]
  wire [2:0] _T_527 = laddr_reg == addrMetaMem_listenAddr_MPORT_3_data ? 3'h4 : {{1'd0}, _T_525}; // @[DFCTableD.scala 72:21]
  wire [2:0] _T_529 = laddr_reg == addrMetaMem_listenAddr_MPORT_4_data ? 3'h5 : _T_527; // @[DFCTableD.scala 72:21]
  wire [2:0] _T_531 = laddr_reg == addrMetaMem_listenAddr_MPORT_5_data ? 3'h6 : _T_529; // @[DFCTableD.scala 72:21]
  wire [2:0] _T_533 = laddr_reg == addrMetaMem_listenAddr_MPORT_6_data ? 3'h7 : _T_531; // @[DFCTableD.scala 72:21]
  wire [3:0] _T_535 = laddr_reg == addrMetaMem_listenAddr_MPORT_7_data ? 4'h8 : {{1'd0}, _T_533}; // @[DFCTableD.scala 72:21]
  wire [3:0] _T_537 = laddr_reg == addrMetaMem_listenAddr_MPORT_8_data ? 4'h9 : _T_535; // @[DFCTableD.scala 72:21]
  wire [3:0] _T_539 = laddr_reg == addrMetaMem_listenAddr_MPORT_9_data ? 4'ha : _T_537; // @[DFCTableD.scala 72:21]
  wire [3:0] _T_541 = laddr_reg == addrMetaMem_listenAddr_MPORT_10_data ? 4'hb : _T_539; // @[DFCTableD.scala 72:21]
  wire [3:0] _T_543 = laddr_reg == addrMetaMem_listenAddr_MPORT_11_data ? 4'hc : _T_541; // @[DFCTableD.scala 72:21]
  wire [3:0] _T_545 = laddr_reg == addrMetaMem_listenAddr_MPORT_12_data ? 4'hd : _T_543; // @[DFCTableD.scala 72:21]
  wire [3:0] _T_547 = laddr_reg == addrMetaMem_listenAddr_MPORT_13_data ? 4'he : _T_545; // @[DFCTableD.scala 72:21]
  wire [3:0] _T_549 = laddr_reg == addrMetaMem_listenAddr_MPORT_14_data ? 4'hf : _T_547; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_551 = laddr_reg == addrMetaMem_listenAddr_MPORT_15_data ? 5'h10 : {{1'd0}, _T_549}; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_553 = laddr_reg == addrMetaMem_listenAddr_MPORT_16_data ? 5'h11 : _T_551; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_555 = laddr_reg == addrMetaMem_listenAddr_MPORT_17_data ? 5'h12 : _T_553; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_557 = laddr_reg == addrMetaMem_listenAddr_MPORT_18_data ? 5'h13 : _T_555; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_559 = laddr_reg == addrMetaMem_listenAddr_MPORT_19_data ? 5'h14 : _T_557; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_561 = laddr_reg == addrMetaMem_listenAddr_MPORT_20_data ? 5'h15 : _T_559; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_563 = laddr_reg == addrMetaMem_listenAddr_MPORT_21_data ? 5'h16 : _T_561; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_565 = laddr_reg == addrMetaMem_listenAddr_MPORT_22_data ? 5'h17 : _T_563; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_567 = laddr_reg == addrMetaMem_listenAddr_MPORT_23_data ? 5'h18 : _T_565; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_569 = laddr_reg == addrMetaMem_listenAddr_MPORT_24_data ? 5'h19 : _T_567; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_571 = laddr_reg == addrMetaMem_listenAddr_MPORT_25_data ? 5'h1a : _T_569; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_573 = laddr_reg == addrMetaMem_listenAddr_MPORT_26_data ? 5'h1b : _T_571; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_575 = laddr_reg == addrMetaMem_listenAddr_MPORT_27_data ? 5'h1c : _T_573; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_577 = laddr_reg == addrMetaMem_listenAddr_MPORT_28_data ? 5'h1d : _T_575; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_579 = laddr_reg == addrMetaMem_listenAddr_MPORT_29_data ? 5'h1e : _T_577; // @[DFCTableD.scala 72:21]
  wire [4:0] _T_581 = laddr_reg == addrMetaMem_listenAddr_MPORT_30_data ? 5'h1f : _T_579; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_583 = laddr_reg == addrMetaMem_listenAddr_MPORT_31_data ? 6'h20 : {{1'd0}, _T_581}; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_585 = laddr_reg == addrMetaMem_listenAddr_MPORT_32_data ? 6'h21 : _T_583; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_587 = laddr_reg == addrMetaMem_listenAddr_MPORT_33_data ? 6'h22 : _T_585; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_589 = laddr_reg == addrMetaMem_listenAddr_MPORT_34_data ? 6'h23 : _T_587; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_591 = laddr_reg == addrMetaMem_listenAddr_MPORT_35_data ? 6'h24 : _T_589; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_593 = laddr_reg == addrMetaMem_listenAddr_MPORT_36_data ? 6'h25 : _T_591; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_595 = laddr_reg == addrMetaMem_listenAddr_MPORT_37_data ? 6'h26 : _T_593; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_597 = laddr_reg == addrMetaMem_listenAddr_MPORT_38_data ? 6'h27 : _T_595; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_599 = laddr_reg == addrMetaMem_listenAddr_MPORT_39_data ? 6'h28 : _T_597; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_601 = laddr_reg == addrMetaMem_listenAddr_MPORT_40_data ? 6'h29 : _T_599; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_603 = laddr_reg == addrMetaMem_listenAddr_MPORT_41_data ? 6'h2a : _T_601; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_605 = laddr_reg == addrMetaMem_listenAddr_MPORT_42_data ? 6'h2b : _T_603; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_607 = laddr_reg == addrMetaMem_listenAddr_MPORT_43_data ? 6'h2c : _T_605; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_609 = laddr_reg == addrMetaMem_listenAddr_MPORT_44_data ? 6'h2d : _T_607; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_611 = laddr_reg == addrMetaMem_listenAddr_MPORT_45_data ? 6'h2e : _T_609; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_613 = laddr_reg == addrMetaMem_listenAddr_MPORT_46_data ? 6'h2f : _T_611; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_615 = laddr_reg == addrMetaMem_listenAddr_MPORT_47_data ? 6'h30 : _T_613; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_617 = laddr_reg == addrMetaMem_listenAddr_MPORT_48_data ? 6'h31 : _T_615; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_619 = laddr_reg == addrMetaMem_listenAddr_MPORT_49_data ? 6'h32 : _T_617; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_621 = laddr_reg == addrMetaMem_listenAddr_MPORT_50_data ? 6'h33 : _T_619; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_623 = laddr_reg == addrMetaMem_listenAddr_MPORT_51_data ? 6'h34 : _T_621; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_625 = laddr_reg == addrMetaMem_listenAddr_MPORT_52_data ? 6'h35 : _T_623; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_627 = laddr_reg == addrMetaMem_listenAddr_MPORT_53_data ? 6'h36 : _T_625; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_629 = laddr_reg == addrMetaMem_listenAddr_MPORT_54_data ? 6'h37 : _T_627; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_631 = laddr_reg == addrMetaMem_listenAddr_MPORT_55_data ? 6'h38 : _T_629; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_633 = laddr_reg == addrMetaMem_listenAddr_MPORT_56_data ? 6'h39 : _T_631; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_635 = laddr_reg == addrMetaMem_listenAddr_MPORT_57_data ? 6'h3a : _T_633; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_637 = laddr_reg == addrMetaMem_listenAddr_MPORT_58_data ? 6'h3b : _T_635; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_639 = laddr_reg == addrMetaMem_listenAddr_MPORT_59_data ? 6'h3c : _T_637; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_641 = laddr_reg == addrMetaMem_listenAddr_MPORT_60_data ? 6'h3d : _T_639; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_643 = laddr_reg == addrMetaMem_listenAddr_MPORT_61_data ? 6'h3e : _T_641; // @[DFCTableD.scala 72:21]
  wire [5:0] _T_645 = laddr_reg == addrMetaMem_listenAddr_MPORT_62_data ? 6'h3f : _T_643; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_647 = laddr_reg == addrMetaMem_listenAddr_MPORT_63_data ? 7'h40 : {{1'd0}, _T_645}; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_649 = laddr_reg == addrMetaMem_listenAddr_MPORT_64_data ? 7'h41 : _T_647; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_651 = laddr_reg == addrMetaMem_listenAddr_MPORT_65_data ? 7'h42 : _T_649; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_653 = laddr_reg == addrMetaMem_listenAddr_MPORT_66_data ? 7'h43 : _T_651; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_655 = laddr_reg == addrMetaMem_listenAddr_MPORT_67_data ? 7'h44 : _T_653; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_657 = laddr_reg == addrMetaMem_listenAddr_MPORT_68_data ? 7'h45 : _T_655; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_659 = laddr_reg == addrMetaMem_listenAddr_MPORT_69_data ? 7'h46 : _T_657; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_661 = laddr_reg == addrMetaMem_listenAddr_MPORT_70_data ? 7'h47 : _T_659; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_663 = laddr_reg == addrMetaMem_listenAddr_MPORT_71_data ? 7'h48 : _T_661; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_665 = laddr_reg == addrMetaMem_listenAddr_MPORT_72_data ? 7'h49 : _T_663; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_667 = laddr_reg == addrMetaMem_listenAddr_MPORT_73_data ? 7'h4a : _T_665; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_669 = laddr_reg == addrMetaMem_listenAddr_MPORT_74_data ? 7'h4b : _T_667; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_671 = laddr_reg == addrMetaMem_listenAddr_MPORT_75_data ? 7'h4c : _T_669; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_673 = laddr_reg == addrMetaMem_listenAddr_MPORT_76_data ? 7'h4d : _T_671; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_675 = laddr_reg == addrMetaMem_listenAddr_MPORT_77_data ? 7'h4e : _T_673; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_677 = laddr_reg == addrMetaMem_listenAddr_MPORT_78_data ? 7'h4f : _T_675; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_679 = laddr_reg == addrMetaMem_listenAddr_MPORT_79_data ? 7'h50 : _T_677; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_681 = laddr_reg == addrMetaMem_listenAddr_MPORT_80_data ? 7'h51 : _T_679; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_683 = laddr_reg == addrMetaMem_listenAddr_MPORT_81_data ? 7'h52 : _T_681; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_685 = laddr_reg == addrMetaMem_listenAddr_MPORT_82_data ? 7'h53 : _T_683; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_687 = laddr_reg == addrMetaMem_listenAddr_MPORT_83_data ? 7'h54 : _T_685; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_689 = laddr_reg == addrMetaMem_listenAddr_MPORT_84_data ? 7'h55 : _T_687; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_691 = laddr_reg == addrMetaMem_listenAddr_MPORT_85_data ? 7'h56 : _T_689; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_693 = laddr_reg == addrMetaMem_listenAddr_MPORT_86_data ? 7'h57 : _T_691; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_695 = laddr_reg == addrMetaMem_listenAddr_MPORT_87_data ? 7'h58 : _T_693; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_697 = laddr_reg == addrMetaMem_listenAddr_MPORT_88_data ? 7'h59 : _T_695; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_699 = laddr_reg == addrMetaMem_listenAddr_MPORT_89_data ? 7'h5a : _T_697; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_701 = laddr_reg == addrMetaMem_listenAddr_MPORT_90_data ? 7'h5b : _T_699; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_703 = laddr_reg == addrMetaMem_listenAddr_MPORT_91_data ? 7'h5c : _T_701; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_705 = laddr_reg == addrMetaMem_listenAddr_MPORT_92_data ? 7'h5d : _T_703; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_707 = laddr_reg == addrMetaMem_listenAddr_MPORT_93_data ? 7'h5e : _T_705; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_709 = laddr_reg == addrMetaMem_listenAddr_MPORT_94_data ? 7'h5f : _T_707; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_711 = laddr_reg == addrMetaMem_listenAddr_MPORT_95_data ? 7'h60 : _T_709; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_713 = laddr_reg == addrMetaMem_listenAddr_MPORT_96_data ? 7'h61 : _T_711; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_715 = laddr_reg == addrMetaMem_listenAddr_MPORT_97_data ? 7'h62 : _T_713; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_717 = laddr_reg == addrMetaMem_listenAddr_MPORT_98_data ? 7'h63 : _T_715; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_719 = laddr_reg == addrMetaMem_listenAddr_MPORT_99_data ? 7'h64 : _T_717; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_721 = laddr_reg == addrMetaMem_listenAddr_MPORT_100_data ? 7'h65 : _T_719; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_723 = laddr_reg == addrMetaMem_listenAddr_MPORT_101_data ? 7'h66 : _T_721; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_725 = laddr_reg == addrMetaMem_listenAddr_MPORT_102_data ? 7'h67 : _T_723; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_727 = laddr_reg == addrMetaMem_listenAddr_MPORT_103_data ? 7'h68 : _T_725; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_729 = laddr_reg == addrMetaMem_listenAddr_MPORT_104_data ? 7'h69 : _T_727; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_731 = laddr_reg == addrMetaMem_listenAddr_MPORT_105_data ? 7'h6a : _T_729; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_733 = laddr_reg == addrMetaMem_listenAddr_MPORT_106_data ? 7'h6b : _T_731; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_735 = laddr_reg == addrMetaMem_listenAddr_MPORT_107_data ? 7'h6c : _T_733; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_737 = laddr_reg == addrMetaMem_listenAddr_MPORT_108_data ? 7'h6d : _T_735; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_739 = laddr_reg == addrMetaMem_listenAddr_MPORT_109_data ? 7'h6e : _T_737; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_741 = laddr_reg == addrMetaMem_listenAddr_MPORT_110_data ? 7'h6f : _T_739; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_743 = laddr_reg == addrMetaMem_listenAddr_MPORT_111_data ? 7'h70 : _T_741; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_745 = laddr_reg == addrMetaMem_listenAddr_MPORT_112_data ? 7'h71 : _T_743; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_747 = laddr_reg == addrMetaMem_listenAddr_MPORT_113_data ? 7'h72 : _T_745; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_749 = laddr_reg == addrMetaMem_listenAddr_MPORT_114_data ? 7'h73 : _T_747; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_751 = laddr_reg == addrMetaMem_listenAddr_MPORT_115_data ? 7'h74 : _T_749; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_753 = laddr_reg == addrMetaMem_listenAddr_MPORT_116_data ? 7'h75 : _T_751; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_755 = laddr_reg == addrMetaMem_listenAddr_MPORT_117_data ? 7'h76 : _T_753; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_757 = laddr_reg == addrMetaMem_listenAddr_MPORT_118_data ? 7'h77 : _T_755; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_759 = laddr_reg == addrMetaMem_listenAddr_MPORT_119_data ? 7'h78 : _T_757; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_761 = laddr_reg == addrMetaMem_listenAddr_MPORT_120_data ? 7'h79 : _T_759; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_763 = laddr_reg == addrMetaMem_listenAddr_MPORT_121_data ? 7'h7a : _T_761; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_765 = laddr_reg == addrMetaMem_listenAddr_MPORT_122_data ? 7'h7b : _T_763; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_767 = laddr_reg == addrMetaMem_listenAddr_MPORT_123_data ? 7'h7c : _T_765; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_769 = laddr_reg == addrMetaMem_listenAddr_MPORT_124_data ? 7'h7d : _T_767; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_771 = laddr_reg == addrMetaMem_listenAddr_MPORT_125_data ? 7'h7e : _T_769; // @[DFCTableD.scala 72:21]
  wire [6:0] _T_773 = laddr_reg == addrMetaMem_listenAddr_MPORT_126_data ? 7'h7f : _T_771; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_775 = laddr_reg == addrMetaMem_listenAddr_MPORT_127_data ? 8'h80 : {{1'd0}, _T_773}; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_777 = laddr_reg == addrMetaMem_listenAddr_MPORT_128_data ? 8'h81 : _T_775; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_779 = laddr_reg == addrMetaMem_listenAddr_MPORT_129_data ? 8'h82 : _T_777; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_781 = laddr_reg == addrMetaMem_listenAddr_MPORT_130_data ? 8'h83 : _T_779; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_783 = laddr_reg == addrMetaMem_listenAddr_MPORT_131_data ? 8'h84 : _T_781; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_785 = laddr_reg == addrMetaMem_listenAddr_MPORT_132_data ? 8'h85 : _T_783; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_787 = laddr_reg == addrMetaMem_listenAddr_MPORT_133_data ? 8'h86 : _T_785; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_789 = laddr_reg == addrMetaMem_listenAddr_MPORT_134_data ? 8'h87 : _T_787; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_791 = laddr_reg == addrMetaMem_listenAddr_MPORT_135_data ? 8'h88 : _T_789; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_793 = laddr_reg == addrMetaMem_listenAddr_MPORT_136_data ? 8'h89 : _T_791; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_795 = laddr_reg == addrMetaMem_listenAddr_MPORT_137_data ? 8'h8a : _T_793; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_797 = laddr_reg == addrMetaMem_listenAddr_MPORT_138_data ? 8'h8b : _T_795; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_799 = laddr_reg == addrMetaMem_listenAddr_MPORT_139_data ? 8'h8c : _T_797; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_801 = laddr_reg == addrMetaMem_listenAddr_MPORT_140_data ? 8'h8d : _T_799; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_803 = laddr_reg == addrMetaMem_listenAddr_MPORT_141_data ? 8'h8e : _T_801; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_805 = laddr_reg == addrMetaMem_listenAddr_MPORT_142_data ? 8'h8f : _T_803; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_807 = laddr_reg == addrMetaMem_listenAddr_MPORT_143_data ? 8'h90 : _T_805; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_809 = laddr_reg == addrMetaMem_listenAddr_MPORT_144_data ? 8'h91 : _T_807; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_811 = laddr_reg == addrMetaMem_listenAddr_MPORT_145_data ? 8'h92 : _T_809; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_813 = laddr_reg == addrMetaMem_listenAddr_MPORT_146_data ? 8'h93 : _T_811; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_815 = laddr_reg == addrMetaMem_listenAddr_MPORT_147_data ? 8'h94 : _T_813; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_817 = laddr_reg == addrMetaMem_listenAddr_MPORT_148_data ? 8'h95 : _T_815; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_819 = laddr_reg == addrMetaMem_listenAddr_MPORT_149_data ? 8'h96 : _T_817; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_821 = laddr_reg == addrMetaMem_listenAddr_MPORT_150_data ? 8'h97 : _T_819; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_823 = laddr_reg == addrMetaMem_listenAddr_MPORT_151_data ? 8'h98 : _T_821; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_825 = laddr_reg == addrMetaMem_listenAddr_MPORT_152_data ? 8'h99 : _T_823; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_827 = laddr_reg == addrMetaMem_listenAddr_MPORT_153_data ? 8'h9a : _T_825; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_829 = laddr_reg == addrMetaMem_listenAddr_MPORT_154_data ? 8'h9b : _T_827; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_831 = laddr_reg == addrMetaMem_listenAddr_MPORT_155_data ? 8'h9c : _T_829; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_833 = laddr_reg == addrMetaMem_listenAddr_MPORT_156_data ? 8'h9d : _T_831; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_835 = laddr_reg == addrMetaMem_listenAddr_MPORT_157_data ? 8'h9e : _T_833; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_837 = laddr_reg == addrMetaMem_listenAddr_MPORT_158_data ? 8'h9f : _T_835; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_839 = laddr_reg == addrMetaMem_listenAddr_MPORT_159_data ? 8'ha0 : _T_837; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_841 = laddr_reg == addrMetaMem_listenAddr_MPORT_160_data ? 8'ha1 : _T_839; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_843 = laddr_reg == addrMetaMem_listenAddr_MPORT_161_data ? 8'ha2 : _T_841; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_845 = laddr_reg == addrMetaMem_listenAddr_MPORT_162_data ? 8'ha3 : _T_843; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_847 = laddr_reg == addrMetaMem_listenAddr_MPORT_163_data ? 8'ha4 : _T_845; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_849 = laddr_reg == addrMetaMem_listenAddr_MPORT_164_data ? 8'ha5 : _T_847; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_851 = laddr_reg == addrMetaMem_listenAddr_MPORT_165_data ? 8'ha6 : _T_849; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_853 = laddr_reg == addrMetaMem_listenAddr_MPORT_166_data ? 8'ha7 : _T_851; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_855 = laddr_reg == addrMetaMem_listenAddr_MPORT_167_data ? 8'ha8 : _T_853; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_857 = laddr_reg == addrMetaMem_listenAddr_MPORT_168_data ? 8'ha9 : _T_855; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_859 = laddr_reg == addrMetaMem_listenAddr_MPORT_169_data ? 8'haa : _T_857; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_861 = laddr_reg == addrMetaMem_listenAddr_MPORT_170_data ? 8'hab : _T_859; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_863 = laddr_reg == addrMetaMem_listenAddr_MPORT_171_data ? 8'hac : _T_861; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_865 = laddr_reg == addrMetaMem_listenAddr_MPORT_172_data ? 8'had : _T_863; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_867 = laddr_reg == addrMetaMem_listenAddr_MPORT_173_data ? 8'hae : _T_865; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_869 = laddr_reg == addrMetaMem_listenAddr_MPORT_174_data ? 8'haf : _T_867; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_871 = laddr_reg == addrMetaMem_listenAddr_MPORT_175_data ? 8'hb0 : _T_869; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_873 = laddr_reg == addrMetaMem_listenAddr_MPORT_176_data ? 8'hb1 : _T_871; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_875 = laddr_reg == addrMetaMem_listenAddr_MPORT_177_data ? 8'hb2 : _T_873; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_877 = laddr_reg == addrMetaMem_listenAddr_MPORT_178_data ? 8'hb3 : _T_875; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_879 = laddr_reg == addrMetaMem_listenAddr_MPORT_179_data ? 8'hb4 : _T_877; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_881 = laddr_reg == addrMetaMem_listenAddr_MPORT_180_data ? 8'hb5 : _T_879; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_883 = laddr_reg == addrMetaMem_listenAddr_MPORT_181_data ? 8'hb6 : _T_881; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_885 = laddr_reg == addrMetaMem_listenAddr_MPORT_182_data ? 8'hb7 : _T_883; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_887 = laddr_reg == addrMetaMem_listenAddr_MPORT_183_data ? 8'hb8 : _T_885; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_889 = laddr_reg == addrMetaMem_listenAddr_MPORT_184_data ? 8'hb9 : _T_887; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_891 = laddr_reg == addrMetaMem_listenAddr_MPORT_185_data ? 8'hba : _T_889; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_893 = laddr_reg == addrMetaMem_listenAddr_MPORT_186_data ? 8'hbb : _T_891; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_895 = laddr_reg == addrMetaMem_listenAddr_MPORT_187_data ? 8'hbc : _T_893; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_897 = laddr_reg == addrMetaMem_listenAddr_MPORT_188_data ? 8'hbd : _T_895; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_899 = laddr_reg == addrMetaMem_listenAddr_MPORT_189_data ? 8'hbe : _T_897; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_901 = laddr_reg == addrMetaMem_listenAddr_MPORT_190_data ? 8'hbf : _T_899; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_903 = laddr_reg == addrMetaMem_listenAddr_MPORT_191_data ? 8'hc0 : _T_901; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_905 = laddr_reg == addrMetaMem_listenAddr_MPORT_192_data ? 8'hc1 : _T_903; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_907 = laddr_reg == addrMetaMem_listenAddr_MPORT_193_data ? 8'hc2 : _T_905; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_909 = laddr_reg == addrMetaMem_listenAddr_MPORT_194_data ? 8'hc3 : _T_907; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_911 = laddr_reg == addrMetaMem_listenAddr_MPORT_195_data ? 8'hc4 : _T_909; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_913 = laddr_reg == addrMetaMem_listenAddr_MPORT_196_data ? 8'hc5 : _T_911; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_915 = laddr_reg == addrMetaMem_listenAddr_MPORT_197_data ? 8'hc6 : _T_913; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_917 = laddr_reg == addrMetaMem_listenAddr_MPORT_198_data ? 8'hc7 : _T_915; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_919 = laddr_reg == addrMetaMem_listenAddr_MPORT_199_data ? 8'hc8 : _T_917; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_921 = laddr_reg == addrMetaMem_listenAddr_MPORT_200_data ? 8'hc9 : _T_919; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_923 = laddr_reg == addrMetaMem_listenAddr_MPORT_201_data ? 8'hca : _T_921; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_925 = laddr_reg == addrMetaMem_listenAddr_MPORT_202_data ? 8'hcb : _T_923; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_927 = laddr_reg == addrMetaMem_listenAddr_MPORT_203_data ? 8'hcc : _T_925; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_929 = laddr_reg == addrMetaMem_listenAddr_MPORT_204_data ? 8'hcd : _T_927; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_931 = laddr_reg == addrMetaMem_listenAddr_MPORT_205_data ? 8'hce : _T_929; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_933 = laddr_reg == addrMetaMem_listenAddr_MPORT_206_data ? 8'hcf : _T_931; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_935 = laddr_reg == addrMetaMem_listenAddr_MPORT_207_data ? 8'hd0 : _T_933; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_937 = laddr_reg == addrMetaMem_listenAddr_MPORT_208_data ? 8'hd1 : _T_935; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_939 = laddr_reg == addrMetaMem_listenAddr_MPORT_209_data ? 8'hd2 : _T_937; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_941 = laddr_reg == addrMetaMem_listenAddr_MPORT_210_data ? 8'hd3 : _T_939; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_943 = laddr_reg == addrMetaMem_listenAddr_MPORT_211_data ? 8'hd4 : _T_941; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_945 = laddr_reg == addrMetaMem_listenAddr_MPORT_212_data ? 8'hd5 : _T_943; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_947 = laddr_reg == addrMetaMem_listenAddr_MPORT_213_data ? 8'hd6 : _T_945; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_949 = laddr_reg == addrMetaMem_listenAddr_MPORT_214_data ? 8'hd7 : _T_947; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_951 = laddr_reg == addrMetaMem_listenAddr_MPORT_215_data ? 8'hd8 : _T_949; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_953 = laddr_reg == addrMetaMem_listenAddr_MPORT_216_data ? 8'hd9 : _T_951; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_955 = laddr_reg == addrMetaMem_listenAddr_MPORT_217_data ? 8'hda : _T_953; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_957 = laddr_reg == addrMetaMem_listenAddr_MPORT_218_data ? 8'hdb : _T_955; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_959 = laddr_reg == addrMetaMem_listenAddr_MPORT_219_data ? 8'hdc : _T_957; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_961 = laddr_reg == addrMetaMem_listenAddr_MPORT_220_data ? 8'hdd : _T_959; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_963 = laddr_reg == addrMetaMem_listenAddr_MPORT_221_data ? 8'hde : _T_961; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_965 = laddr_reg == addrMetaMem_listenAddr_MPORT_222_data ? 8'hdf : _T_963; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_967 = laddr_reg == addrMetaMem_listenAddr_MPORT_223_data ? 8'he0 : _T_965; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_969 = laddr_reg == addrMetaMem_listenAddr_MPORT_224_data ? 8'he1 : _T_967; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_971 = laddr_reg == addrMetaMem_listenAddr_MPORT_225_data ? 8'he2 : _T_969; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_973 = laddr_reg == addrMetaMem_listenAddr_MPORT_226_data ? 8'he3 : _T_971; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_975 = laddr_reg == addrMetaMem_listenAddr_MPORT_227_data ? 8'he4 : _T_973; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_977 = laddr_reg == addrMetaMem_listenAddr_MPORT_228_data ? 8'he5 : _T_975; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_979 = laddr_reg == addrMetaMem_listenAddr_MPORT_229_data ? 8'he6 : _T_977; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_981 = laddr_reg == addrMetaMem_listenAddr_MPORT_230_data ? 8'he7 : _T_979; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_983 = laddr_reg == addrMetaMem_listenAddr_MPORT_231_data ? 8'he8 : _T_981; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_985 = laddr_reg == addrMetaMem_listenAddr_MPORT_232_data ? 8'he9 : _T_983; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_987 = laddr_reg == addrMetaMem_listenAddr_MPORT_233_data ? 8'hea : _T_985; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_989 = laddr_reg == addrMetaMem_listenAddr_MPORT_234_data ? 8'heb : _T_987; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_991 = laddr_reg == addrMetaMem_listenAddr_MPORT_235_data ? 8'hec : _T_989; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_993 = laddr_reg == addrMetaMem_listenAddr_MPORT_236_data ? 8'hed : _T_991; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_995 = laddr_reg == addrMetaMem_listenAddr_MPORT_237_data ? 8'hee : _T_993; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_997 = laddr_reg == addrMetaMem_listenAddr_MPORT_238_data ? 8'hef : _T_995; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_999 = laddr_reg == addrMetaMem_listenAddr_MPORT_239_data ? 8'hf0 : _T_997; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_1001 = laddr_reg == addrMetaMem_listenAddr_MPORT_240_data ? 8'hf1 : _T_999; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_1003 = laddr_reg == addrMetaMem_listenAddr_MPORT_241_data ? 8'hf2 : _T_1001; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_1005 = laddr_reg == addrMetaMem_listenAddr_MPORT_242_data ? 8'hf3 : _T_1003; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_1007 = laddr_reg == addrMetaMem_listenAddr_MPORT_243_data ? 8'hf4 : _T_1005; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_1009 = laddr_reg == addrMetaMem_listenAddr_MPORT_244_data ? 8'hf5 : _T_1007; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_1011 = laddr_reg == addrMetaMem_listenAddr_MPORT_245_data ? 8'hf6 : _T_1009; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_1013 = laddr_reg == addrMetaMem_listenAddr_MPORT_246_data ? 8'hf7 : _T_1011; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_1015 = laddr_reg == addrMetaMem_listenAddr_MPORT_247_data ? 8'hf8 : _T_1013; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_1017 = laddr_reg == addrMetaMem_listenAddr_MPORT_248_data ? 8'hf9 : _T_1015; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_1019 = laddr_reg == addrMetaMem_listenAddr_MPORT_249_data ? 8'hfa : _T_1017; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_1021 = laddr_reg == addrMetaMem_listenAddr_MPORT_250_data ? 8'hfb : _T_1019; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_1023 = laddr_reg == addrMetaMem_listenAddr_MPORT_251_data ? 8'hfc : _T_1021; // @[DFCTableD.scala 72:21]
  wire [7:0] _T_1025 = laddr_reg == addrMetaMem_listenAddr_MPORT_252_data ? 8'hfd : _T_1023; // @[DFCTableD.scala 72:21]
  wire  _T_1028 = laddr_reg == addrMetaMem_listenAddr_MPORT_254_data; // @[DFCTableD.scala 72:32]
  wire [255:0] _T_1031 = tableD_valid >> match_Id; // @[DFCTableD.scala 77:53]
  wire  notMatched = match_Id == 8'h0 | ~_T_1031[0]; // @[DFCTableD.scala 77:37]
  wire  _T_1034 = state == 3'h1; // @[DFCTableD.scala 89:14]
  wire [255:0] _T_1035 = 256'h1 << tableD_Id; // @[DFCTableD.scala 92:40]
  wire [255:0] _T_1036 = tableD_valid | _T_1035; // @[DFCTableD.scala 92:40]
  wire [255:0] _T_1037 = ~tableD_valid; // @[DFCTableD.scala 92:40]
  wire  _T_1042 = ~reset; // @[DFCTableD.scala 93:11]
  wire  _T_1046 = laststate != 3'h5; // @[DFCTableD.scala 96:40]
  wire  _T_1047 = _T & laststate != 3'h5; // @[DFCTableD.scala 96:27]
  wire [255:0] _T_1048 = 256'h1 << match_Id; // @[DFCTableD.scala 99:40]
  wire [255:0] _T_1051 = _T_1037 | _T_1048; // @[DFCTableD.scala 99:40]
  wire [255:0] _T_1052 = ~_T_1051; // @[DFCTableD.scala 99:40]
  wire  _T_1058 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1059 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_1060 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_1061 = io_tableA_wresp_ready & io_tableA_wresp_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_22 = _T_1061 ? 3'h0 : state; // @[DFCTableD.scala 121:35 DFCTableD.scala 122:15 DFCTableD.scala 30:22]
  wire  _T_1062 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_1063 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_1064 = io_tableA_lresp_ready & io_tableA_lresp_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_23 = _T_1064 ? 3'h0 : state; // @[DFCTableD.scala 133:37 DFCTableD.scala 134:17 DFCTableD.scala 30:22]
  wire [2:0] _GEN_26 = notMatched ? _GEN_23 : 3'h5; // @[DFCTableD.scala 130:23 DFCTableD.scala 137:15]
  wire  _T_1065 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_27 = _T_1064 ? 3'h3 : state; // @[DFCTableD.scala 143:35 DFCTableD.scala 144:15 DFCTableD.scala 30:22]
  wire  _GEN_29 = _T_1065 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67 DFCTableD.scala 142:35 DFCTableD.scala 51:31]
  wire [2:0] _GEN_30 = _T_1065 ? _GEN_27 : state; // @[Conditional.scala 39:67 DFCTableD.scala 30:22]
  wire  _GEN_31 = _T_1063 ? notMatched : _T_1065; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_33 = _T_1063 ? _GEN_26 : _GEN_30; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_34 = _T_1062 ? 3'h4 : _GEN_33; // @[Conditional.scala 39:67 DFCTableD.scala 127:13]
  wire  _GEN_35 = _T_1062 ? 1'h0 : _GEN_31; // @[Conditional.scala 39:67 DFCTableD.scala 50:25]
  wire  _GEN_40 = _T_1060 ? 1'h0 : _GEN_35; // @[Conditional.scala 39:67 DFCTableD.scala 50:25]
  wire  _GEN_43 = _T_1059 ? 1'h0 : _T_1060; // @[Conditional.scala 39:67 DFCTableD.scala 47:25]
  wire  _GEN_44 = _T_1059 ? 1'h0 : _T_1060 & notEmpty; // @[Conditional.scala 39:67 DFCTableD.scala 48:25]
  wire  _GEN_45 = _T_1059 ? 1'h0 : _GEN_40; // @[Conditional.scala 39:67 DFCTableD.scala 50:25]
  wire  _GEN_46 = _T_1059 | (_T_1060 | (_T_1062 | (_T_1063 | _GEN_29))); // @[Conditional.scala 39:67 DFCTableD.scala 51:31]
  assign addrMetaMem_listenAddr_MPORT_addr = 8'h1;
  assign addrMetaMem_listenAddr_MPORT_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_1_addr = 8'h2;
  assign addrMetaMem_listenAddr_MPORT_1_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_1_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_2_addr = 8'h3;
  assign addrMetaMem_listenAddr_MPORT_2_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_2_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_3_addr = 8'h4;
  assign addrMetaMem_listenAddr_MPORT_3_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_3_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_4_addr = 8'h5;
  assign addrMetaMem_listenAddr_MPORT_4_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_4_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_5_addr = 8'h6;
  assign addrMetaMem_listenAddr_MPORT_5_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_5_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_6_addr = 8'h7;
  assign addrMetaMem_listenAddr_MPORT_6_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_6_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_7_addr = 8'h8;
  assign addrMetaMem_listenAddr_MPORT_7_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_7_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_8_addr = 8'h9;
  assign addrMetaMem_listenAddr_MPORT_8_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_8_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_9_addr = 8'ha;
  assign addrMetaMem_listenAddr_MPORT_9_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_9_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_10_addr = 8'hb;
  assign addrMetaMem_listenAddr_MPORT_10_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_10_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_11_addr = 8'hc;
  assign addrMetaMem_listenAddr_MPORT_11_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_11_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_12_addr = 8'hd;
  assign addrMetaMem_listenAddr_MPORT_12_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_12_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_13_addr = 8'he;
  assign addrMetaMem_listenAddr_MPORT_13_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_13_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_14_addr = 8'hf;
  assign addrMetaMem_listenAddr_MPORT_14_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_14_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_15_addr = 8'h10;
  assign addrMetaMem_listenAddr_MPORT_15_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_15_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_16_addr = 8'h11;
  assign addrMetaMem_listenAddr_MPORT_16_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_16_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_17_addr = 8'h12;
  assign addrMetaMem_listenAddr_MPORT_17_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_17_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_18_addr = 8'h13;
  assign addrMetaMem_listenAddr_MPORT_18_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_18_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_19_addr = 8'h14;
  assign addrMetaMem_listenAddr_MPORT_19_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_19_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_20_addr = 8'h15;
  assign addrMetaMem_listenAddr_MPORT_20_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_20_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_21_addr = 8'h16;
  assign addrMetaMem_listenAddr_MPORT_21_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_21_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_22_addr = 8'h17;
  assign addrMetaMem_listenAddr_MPORT_22_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_22_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_23_addr = 8'h18;
  assign addrMetaMem_listenAddr_MPORT_23_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_23_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_24_addr = 8'h19;
  assign addrMetaMem_listenAddr_MPORT_24_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_24_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_25_addr = 8'h1a;
  assign addrMetaMem_listenAddr_MPORT_25_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_25_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_26_addr = 8'h1b;
  assign addrMetaMem_listenAddr_MPORT_26_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_26_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_27_addr = 8'h1c;
  assign addrMetaMem_listenAddr_MPORT_27_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_27_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_28_addr = 8'h1d;
  assign addrMetaMem_listenAddr_MPORT_28_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_28_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_29_addr = 8'h1e;
  assign addrMetaMem_listenAddr_MPORT_29_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_29_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_30_addr = 8'h1f;
  assign addrMetaMem_listenAddr_MPORT_30_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_30_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_31_addr = 8'h20;
  assign addrMetaMem_listenAddr_MPORT_31_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_31_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_32_addr = 8'h21;
  assign addrMetaMem_listenAddr_MPORT_32_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_32_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_33_addr = 8'h22;
  assign addrMetaMem_listenAddr_MPORT_33_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_33_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_34_addr = 8'h23;
  assign addrMetaMem_listenAddr_MPORT_34_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_34_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_35_addr = 8'h24;
  assign addrMetaMem_listenAddr_MPORT_35_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_35_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_36_addr = 8'h25;
  assign addrMetaMem_listenAddr_MPORT_36_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_36_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_37_addr = 8'h26;
  assign addrMetaMem_listenAddr_MPORT_37_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_37_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_38_addr = 8'h27;
  assign addrMetaMem_listenAddr_MPORT_38_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_38_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_39_addr = 8'h28;
  assign addrMetaMem_listenAddr_MPORT_39_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_39_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_40_addr = 8'h29;
  assign addrMetaMem_listenAddr_MPORT_40_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_40_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_41_addr = 8'h2a;
  assign addrMetaMem_listenAddr_MPORT_41_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_41_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_42_addr = 8'h2b;
  assign addrMetaMem_listenAddr_MPORT_42_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_42_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_43_addr = 8'h2c;
  assign addrMetaMem_listenAddr_MPORT_43_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_43_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_44_addr = 8'h2d;
  assign addrMetaMem_listenAddr_MPORT_44_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_44_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_45_addr = 8'h2e;
  assign addrMetaMem_listenAddr_MPORT_45_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_45_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_46_addr = 8'h2f;
  assign addrMetaMem_listenAddr_MPORT_46_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_46_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_47_addr = 8'h30;
  assign addrMetaMem_listenAddr_MPORT_47_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_47_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_48_addr = 8'h31;
  assign addrMetaMem_listenAddr_MPORT_48_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_48_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_49_addr = 8'h32;
  assign addrMetaMem_listenAddr_MPORT_49_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_49_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_50_addr = 8'h33;
  assign addrMetaMem_listenAddr_MPORT_50_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_50_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_51_addr = 8'h34;
  assign addrMetaMem_listenAddr_MPORT_51_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_51_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_52_addr = 8'h35;
  assign addrMetaMem_listenAddr_MPORT_52_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_52_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_53_addr = 8'h36;
  assign addrMetaMem_listenAddr_MPORT_53_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_53_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_54_addr = 8'h37;
  assign addrMetaMem_listenAddr_MPORT_54_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_54_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_55_addr = 8'h38;
  assign addrMetaMem_listenAddr_MPORT_55_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_55_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_56_addr = 8'h39;
  assign addrMetaMem_listenAddr_MPORT_56_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_56_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_57_addr = 8'h3a;
  assign addrMetaMem_listenAddr_MPORT_57_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_57_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_58_addr = 8'h3b;
  assign addrMetaMem_listenAddr_MPORT_58_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_58_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_59_addr = 8'h3c;
  assign addrMetaMem_listenAddr_MPORT_59_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_59_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_60_addr = 8'h3d;
  assign addrMetaMem_listenAddr_MPORT_60_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_60_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_61_addr = 8'h3e;
  assign addrMetaMem_listenAddr_MPORT_61_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_61_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_62_addr = 8'h3f;
  assign addrMetaMem_listenAddr_MPORT_62_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_62_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_63_addr = 8'h40;
  assign addrMetaMem_listenAddr_MPORT_63_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_63_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_64_addr = 8'h41;
  assign addrMetaMem_listenAddr_MPORT_64_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_64_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_65_addr = 8'h42;
  assign addrMetaMem_listenAddr_MPORT_65_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_65_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_66_addr = 8'h43;
  assign addrMetaMem_listenAddr_MPORT_66_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_66_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_67_addr = 8'h44;
  assign addrMetaMem_listenAddr_MPORT_67_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_67_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_68_addr = 8'h45;
  assign addrMetaMem_listenAddr_MPORT_68_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_68_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_69_addr = 8'h46;
  assign addrMetaMem_listenAddr_MPORT_69_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_69_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_70_addr = 8'h47;
  assign addrMetaMem_listenAddr_MPORT_70_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_70_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_71_addr = 8'h48;
  assign addrMetaMem_listenAddr_MPORT_71_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_71_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_72_addr = 8'h49;
  assign addrMetaMem_listenAddr_MPORT_72_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_72_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_73_addr = 8'h4a;
  assign addrMetaMem_listenAddr_MPORT_73_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_73_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_74_addr = 8'h4b;
  assign addrMetaMem_listenAddr_MPORT_74_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_74_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_75_addr = 8'h4c;
  assign addrMetaMem_listenAddr_MPORT_75_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_75_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_76_addr = 8'h4d;
  assign addrMetaMem_listenAddr_MPORT_76_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_76_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_77_addr = 8'h4e;
  assign addrMetaMem_listenAddr_MPORT_77_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_77_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_78_addr = 8'h4f;
  assign addrMetaMem_listenAddr_MPORT_78_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_78_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_79_addr = 8'h50;
  assign addrMetaMem_listenAddr_MPORT_79_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_79_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_80_addr = 8'h51;
  assign addrMetaMem_listenAddr_MPORT_80_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_80_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_81_addr = 8'h52;
  assign addrMetaMem_listenAddr_MPORT_81_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_81_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_82_addr = 8'h53;
  assign addrMetaMem_listenAddr_MPORT_82_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_82_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_83_addr = 8'h54;
  assign addrMetaMem_listenAddr_MPORT_83_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_83_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_84_addr = 8'h55;
  assign addrMetaMem_listenAddr_MPORT_84_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_84_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_85_addr = 8'h56;
  assign addrMetaMem_listenAddr_MPORT_85_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_85_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_86_addr = 8'h57;
  assign addrMetaMem_listenAddr_MPORT_86_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_86_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_87_addr = 8'h58;
  assign addrMetaMem_listenAddr_MPORT_87_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_87_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_88_addr = 8'h59;
  assign addrMetaMem_listenAddr_MPORT_88_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_88_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_89_addr = 8'h5a;
  assign addrMetaMem_listenAddr_MPORT_89_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_89_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_90_addr = 8'h5b;
  assign addrMetaMem_listenAddr_MPORT_90_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_90_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_91_addr = 8'h5c;
  assign addrMetaMem_listenAddr_MPORT_91_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_91_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_92_addr = 8'h5d;
  assign addrMetaMem_listenAddr_MPORT_92_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_92_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_93_addr = 8'h5e;
  assign addrMetaMem_listenAddr_MPORT_93_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_93_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_94_addr = 8'h5f;
  assign addrMetaMem_listenAddr_MPORT_94_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_94_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_95_addr = 8'h60;
  assign addrMetaMem_listenAddr_MPORT_95_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_95_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_96_addr = 8'h61;
  assign addrMetaMem_listenAddr_MPORT_96_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_96_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_97_addr = 8'h62;
  assign addrMetaMem_listenAddr_MPORT_97_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_97_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_98_addr = 8'h63;
  assign addrMetaMem_listenAddr_MPORT_98_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_98_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_99_addr = 8'h64;
  assign addrMetaMem_listenAddr_MPORT_99_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_99_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_100_addr = 8'h65;
  assign addrMetaMem_listenAddr_MPORT_100_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_100_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_101_addr = 8'h66;
  assign addrMetaMem_listenAddr_MPORT_101_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_101_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_102_addr = 8'h67;
  assign addrMetaMem_listenAddr_MPORT_102_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_102_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_103_addr = 8'h68;
  assign addrMetaMem_listenAddr_MPORT_103_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_103_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_104_addr = 8'h69;
  assign addrMetaMem_listenAddr_MPORT_104_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_104_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_105_addr = 8'h6a;
  assign addrMetaMem_listenAddr_MPORT_105_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_105_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_106_addr = 8'h6b;
  assign addrMetaMem_listenAddr_MPORT_106_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_106_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_107_addr = 8'h6c;
  assign addrMetaMem_listenAddr_MPORT_107_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_107_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_108_addr = 8'h6d;
  assign addrMetaMem_listenAddr_MPORT_108_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_108_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_109_addr = 8'h6e;
  assign addrMetaMem_listenAddr_MPORT_109_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_109_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_110_addr = 8'h6f;
  assign addrMetaMem_listenAddr_MPORT_110_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_110_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_111_addr = 8'h70;
  assign addrMetaMem_listenAddr_MPORT_111_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_111_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_112_addr = 8'h71;
  assign addrMetaMem_listenAddr_MPORT_112_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_112_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_113_addr = 8'h72;
  assign addrMetaMem_listenAddr_MPORT_113_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_113_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_114_addr = 8'h73;
  assign addrMetaMem_listenAddr_MPORT_114_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_114_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_115_addr = 8'h74;
  assign addrMetaMem_listenAddr_MPORT_115_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_115_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_116_addr = 8'h75;
  assign addrMetaMem_listenAddr_MPORT_116_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_116_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_117_addr = 8'h76;
  assign addrMetaMem_listenAddr_MPORT_117_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_117_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_118_addr = 8'h77;
  assign addrMetaMem_listenAddr_MPORT_118_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_118_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_119_addr = 8'h78;
  assign addrMetaMem_listenAddr_MPORT_119_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_119_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_120_addr = 8'h79;
  assign addrMetaMem_listenAddr_MPORT_120_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_120_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_121_addr = 8'h7a;
  assign addrMetaMem_listenAddr_MPORT_121_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_121_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_122_addr = 8'h7b;
  assign addrMetaMem_listenAddr_MPORT_122_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_122_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_123_addr = 8'h7c;
  assign addrMetaMem_listenAddr_MPORT_123_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_123_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_124_addr = 8'h7d;
  assign addrMetaMem_listenAddr_MPORT_124_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_124_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_125_addr = 8'h7e;
  assign addrMetaMem_listenAddr_MPORT_125_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_125_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_126_addr = 8'h7f;
  assign addrMetaMem_listenAddr_MPORT_126_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_126_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_127_addr = 8'h80;
  assign addrMetaMem_listenAddr_MPORT_127_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_127_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_128_addr = 8'h81;
  assign addrMetaMem_listenAddr_MPORT_128_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_128_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_129_addr = 8'h82;
  assign addrMetaMem_listenAddr_MPORT_129_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_129_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_130_addr = 8'h83;
  assign addrMetaMem_listenAddr_MPORT_130_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_130_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_131_addr = 8'h84;
  assign addrMetaMem_listenAddr_MPORT_131_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_131_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_132_addr = 8'h85;
  assign addrMetaMem_listenAddr_MPORT_132_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_132_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_133_addr = 8'h86;
  assign addrMetaMem_listenAddr_MPORT_133_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_133_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_134_addr = 8'h87;
  assign addrMetaMem_listenAddr_MPORT_134_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_134_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_135_addr = 8'h88;
  assign addrMetaMem_listenAddr_MPORT_135_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_135_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_136_addr = 8'h89;
  assign addrMetaMem_listenAddr_MPORT_136_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_136_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_137_addr = 8'h8a;
  assign addrMetaMem_listenAddr_MPORT_137_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_137_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_138_addr = 8'h8b;
  assign addrMetaMem_listenAddr_MPORT_138_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_138_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_139_addr = 8'h8c;
  assign addrMetaMem_listenAddr_MPORT_139_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_139_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_140_addr = 8'h8d;
  assign addrMetaMem_listenAddr_MPORT_140_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_140_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_141_addr = 8'h8e;
  assign addrMetaMem_listenAddr_MPORT_141_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_141_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_142_addr = 8'h8f;
  assign addrMetaMem_listenAddr_MPORT_142_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_142_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_143_addr = 8'h90;
  assign addrMetaMem_listenAddr_MPORT_143_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_143_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_144_addr = 8'h91;
  assign addrMetaMem_listenAddr_MPORT_144_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_144_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_145_addr = 8'h92;
  assign addrMetaMem_listenAddr_MPORT_145_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_145_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_146_addr = 8'h93;
  assign addrMetaMem_listenAddr_MPORT_146_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_146_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_147_addr = 8'h94;
  assign addrMetaMem_listenAddr_MPORT_147_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_147_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_148_addr = 8'h95;
  assign addrMetaMem_listenAddr_MPORT_148_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_148_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_149_addr = 8'h96;
  assign addrMetaMem_listenAddr_MPORT_149_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_149_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_150_addr = 8'h97;
  assign addrMetaMem_listenAddr_MPORT_150_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_150_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_151_addr = 8'h98;
  assign addrMetaMem_listenAddr_MPORT_151_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_151_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_152_addr = 8'h99;
  assign addrMetaMem_listenAddr_MPORT_152_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_152_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_153_addr = 8'h9a;
  assign addrMetaMem_listenAddr_MPORT_153_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_153_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_154_addr = 8'h9b;
  assign addrMetaMem_listenAddr_MPORT_154_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_154_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_155_addr = 8'h9c;
  assign addrMetaMem_listenAddr_MPORT_155_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_155_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_156_addr = 8'h9d;
  assign addrMetaMem_listenAddr_MPORT_156_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_156_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_157_addr = 8'h9e;
  assign addrMetaMem_listenAddr_MPORT_157_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_157_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_158_addr = 8'h9f;
  assign addrMetaMem_listenAddr_MPORT_158_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_158_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_159_addr = 8'ha0;
  assign addrMetaMem_listenAddr_MPORT_159_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_159_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_160_addr = 8'ha1;
  assign addrMetaMem_listenAddr_MPORT_160_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_160_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_161_addr = 8'ha2;
  assign addrMetaMem_listenAddr_MPORT_161_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_161_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_162_addr = 8'ha3;
  assign addrMetaMem_listenAddr_MPORT_162_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_162_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_163_addr = 8'ha4;
  assign addrMetaMem_listenAddr_MPORT_163_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_163_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_164_addr = 8'ha5;
  assign addrMetaMem_listenAddr_MPORT_164_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_164_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_165_addr = 8'ha6;
  assign addrMetaMem_listenAddr_MPORT_165_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_165_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_166_addr = 8'ha7;
  assign addrMetaMem_listenAddr_MPORT_166_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_166_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_167_addr = 8'ha8;
  assign addrMetaMem_listenAddr_MPORT_167_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_167_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_168_addr = 8'ha9;
  assign addrMetaMem_listenAddr_MPORT_168_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_168_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_169_addr = 8'haa;
  assign addrMetaMem_listenAddr_MPORT_169_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_169_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_170_addr = 8'hab;
  assign addrMetaMem_listenAddr_MPORT_170_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_170_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_171_addr = 8'hac;
  assign addrMetaMem_listenAddr_MPORT_171_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_171_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_172_addr = 8'had;
  assign addrMetaMem_listenAddr_MPORT_172_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_172_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_173_addr = 8'hae;
  assign addrMetaMem_listenAddr_MPORT_173_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_173_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_174_addr = 8'haf;
  assign addrMetaMem_listenAddr_MPORT_174_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_174_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_175_addr = 8'hb0;
  assign addrMetaMem_listenAddr_MPORT_175_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_175_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_176_addr = 8'hb1;
  assign addrMetaMem_listenAddr_MPORT_176_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_176_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_177_addr = 8'hb2;
  assign addrMetaMem_listenAddr_MPORT_177_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_177_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_178_addr = 8'hb3;
  assign addrMetaMem_listenAddr_MPORT_178_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_178_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_179_addr = 8'hb4;
  assign addrMetaMem_listenAddr_MPORT_179_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_179_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_180_addr = 8'hb5;
  assign addrMetaMem_listenAddr_MPORT_180_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_180_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_181_addr = 8'hb6;
  assign addrMetaMem_listenAddr_MPORT_181_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_181_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_182_addr = 8'hb7;
  assign addrMetaMem_listenAddr_MPORT_182_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_182_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_183_addr = 8'hb8;
  assign addrMetaMem_listenAddr_MPORT_183_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_183_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_184_addr = 8'hb9;
  assign addrMetaMem_listenAddr_MPORT_184_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_184_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_185_addr = 8'hba;
  assign addrMetaMem_listenAddr_MPORT_185_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_185_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_186_addr = 8'hbb;
  assign addrMetaMem_listenAddr_MPORT_186_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_186_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_187_addr = 8'hbc;
  assign addrMetaMem_listenAddr_MPORT_187_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_187_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_188_addr = 8'hbd;
  assign addrMetaMem_listenAddr_MPORT_188_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_188_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_189_addr = 8'hbe;
  assign addrMetaMem_listenAddr_MPORT_189_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_189_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_190_addr = 8'hbf;
  assign addrMetaMem_listenAddr_MPORT_190_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_190_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_191_addr = 8'hc0;
  assign addrMetaMem_listenAddr_MPORT_191_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_191_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_192_addr = 8'hc1;
  assign addrMetaMem_listenAddr_MPORT_192_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_192_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_193_addr = 8'hc2;
  assign addrMetaMem_listenAddr_MPORT_193_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_193_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_194_addr = 8'hc3;
  assign addrMetaMem_listenAddr_MPORT_194_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_194_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_195_addr = 8'hc4;
  assign addrMetaMem_listenAddr_MPORT_195_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_195_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_196_addr = 8'hc5;
  assign addrMetaMem_listenAddr_MPORT_196_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_196_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_197_addr = 8'hc6;
  assign addrMetaMem_listenAddr_MPORT_197_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_197_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_198_addr = 8'hc7;
  assign addrMetaMem_listenAddr_MPORT_198_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_198_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_199_addr = 8'hc8;
  assign addrMetaMem_listenAddr_MPORT_199_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_199_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_200_addr = 8'hc9;
  assign addrMetaMem_listenAddr_MPORT_200_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_200_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_201_addr = 8'hca;
  assign addrMetaMem_listenAddr_MPORT_201_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_201_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_202_addr = 8'hcb;
  assign addrMetaMem_listenAddr_MPORT_202_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_202_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_203_addr = 8'hcc;
  assign addrMetaMem_listenAddr_MPORT_203_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_203_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_204_addr = 8'hcd;
  assign addrMetaMem_listenAddr_MPORT_204_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_204_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_205_addr = 8'hce;
  assign addrMetaMem_listenAddr_MPORT_205_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_205_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_206_addr = 8'hcf;
  assign addrMetaMem_listenAddr_MPORT_206_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_206_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_207_addr = 8'hd0;
  assign addrMetaMem_listenAddr_MPORT_207_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_207_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_208_addr = 8'hd1;
  assign addrMetaMem_listenAddr_MPORT_208_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_208_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_209_addr = 8'hd2;
  assign addrMetaMem_listenAddr_MPORT_209_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_209_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_210_addr = 8'hd3;
  assign addrMetaMem_listenAddr_MPORT_210_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_210_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_211_addr = 8'hd4;
  assign addrMetaMem_listenAddr_MPORT_211_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_211_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_212_addr = 8'hd5;
  assign addrMetaMem_listenAddr_MPORT_212_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_212_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_213_addr = 8'hd6;
  assign addrMetaMem_listenAddr_MPORT_213_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_213_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_214_addr = 8'hd7;
  assign addrMetaMem_listenAddr_MPORT_214_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_214_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_215_addr = 8'hd8;
  assign addrMetaMem_listenAddr_MPORT_215_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_215_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_216_addr = 8'hd9;
  assign addrMetaMem_listenAddr_MPORT_216_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_216_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_217_addr = 8'hda;
  assign addrMetaMem_listenAddr_MPORT_217_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_217_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_218_addr = 8'hdb;
  assign addrMetaMem_listenAddr_MPORT_218_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_218_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_219_addr = 8'hdc;
  assign addrMetaMem_listenAddr_MPORT_219_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_219_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_220_addr = 8'hdd;
  assign addrMetaMem_listenAddr_MPORT_220_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_220_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_221_addr = 8'hde;
  assign addrMetaMem_listenAddr_MPORT_221_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_221_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_222_addr = 8'hdf;
  assign addrMetaMem_listenAddr_MPORT_222_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_222_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_223_addr = 8'he0;
  assign addrMetaMem_listenAddr_MPORT_223_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_223_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_224_addr = 8'he1;
  assign addrMetaMem_listenAddr_MPORT_224_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_224_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_225_addr = 8'he2;
  assign addrMetaMem_listenAddr_MPORT_225_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_225_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_226_addr = 8'he3;
  assign addrMetaMem_listenAddr_MPORT_226_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_226_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_227_addr = 8'he4;
  assign addrMetaMem_listenAddr_MPORT_227_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_227_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_228_addr = 8'he5;
  assign addrMetaMem_listenAddr_MPORT_228_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_228_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_229_addr = 8'he6;
  assign addrMetaMem_listenAddr_MPORT_229_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_229_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_230_addr = 8'he7;
  assign addrMetaMem_listenAddr_MPORT_230_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_230_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_231_addr = 8'he8;
  assign addrMetaMem_listenAddr_MPORT_231_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_231_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_232_addr = 8'he9;
  assign addrMetaMem_listenAddr_MPORT_232_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_232_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_233_addr = 8'hea;
  assign addrMetaMem_listenAddr_MPORT_233_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_233_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_234_addr = 8'heb;
  assign addrMetaMem_listenAddr_MPORT_234_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_234_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_235_addr = 8'hec;
  assign addrMetaMem_listenAddr_MPORT_235_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_235_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_236_addr = 8'hed;
  assign addrMetaMem_listenAddr_MPORT_236_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_236_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_237_addr = 8'hee;
  assign addrMetaMem_listenAddr_MPORT_237_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_237_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_238_addr = 8'hef;
  assign addrMetaMem_listenAddr_MPORT_238_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_238_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_239_addr = 8'hf0;
  assign addrMetaMem_listenAddr_MPORT_239_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_239_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_240_addr = 8'hf1;
  assign addrMetaMem_listenAddr_MPORT_240_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_240_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_241_addr = 8'hf2;
  assign addrMetaMem_listenAddr_MPORT_241_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_241_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_242_addr = 8'hf3;
  assign addrMetaMem_listenAddr_MPORT_242_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_242_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_243_addr = 8'hf4;
  assign addrMetaMem_listenAddr_MPORT_243_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_243_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_244_addr = 8'hf5;
  assign addrMetaMem_listenAddr_MPORT_244_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_244_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_245_addr = 8'hf6;
  assign addrMetaMem_listenAddr_MPORT_245_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_245_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_246_addr = 8'hf7;
  assign addrMetaMem_listenAddr_MPORT_246_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_246_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_247_addr = 8'hf8;
  assign addrMetaMem_listenAddr_MPORT_247_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_247_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_248_addr = 8'hf9;
  assign addrMetaMem_listenAddr_MPORT_248_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_248_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_249_addr = 8'hfa;
  assign addrMetaMem_listenAddr_MPORT_249_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_249_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_250_addr = 8'hfb;
  assign addrMetaMem_listenAddr_MPORT_250_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_250_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_251_addr = 8'hfc;
  assign addrMetaMem_listenAddr_MPORT_251_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_251_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_252_addr = 8'hfd;
  assign addrMetaMem_listenAddr_MPORT_252_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_252_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_253_addr = 8'hfe;
  assign addrMetaMem_listenAddr_MPORT_253_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_253_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_254_addr = 8'hff;
  assign addrMetaMem_listenAddr_MPORT_254_data = addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_254_addr]; // @[DFCTableD.scala 25:32]
  assign addrMetaMem_listenAddr_MPORT_256_data = laddr_reg;
  assign addrMetaMem_listenAddr_MPORT_256_addr = tableD_Id;
  assign addrMetaMem_listenAddr_MPORT_256_mask = 1'h1;
  assign addrMetaMem_listenAddr_MPORT_256_en = state == 3'h1;
  assign addrMetaMem_listenAddr_MPORT_258_data = 32'h0;
  assign addrMetaMem_listenAddr_MPORT_258_addr = match_Id;
  assign addrMetaMem_listenAddr_MPORT_258_mask = 1'h1;
  assign addrMetaMem_listenAddr_MPORT_258_en = _T & _T_1046;
  assign infoMetaMem_tableAid_MPORT_255_addr = infoMetaMem_tableAid_MPORT_255_addr_pipe_0;
  assign infoMetaMem_tableAid_MPORT_255_data = infoMetaMem_tableAid[infoMetaMem_tableAid_MPORT_255_addr]; // @[DFCTableD.scala 26:32]
  assign infoMetaMem_tableAid_MPORT_257_data = tableAid_reg;
  assign infoMetaMem_tableAid_MPORT_257_addr = tableD_Id;
  assign infoMetaMem_tableAid_MPORT_257_mask = 1'h1;
  assign infoMetaMem_tableAid_MPORT_257_en = state == 3'h1;
  assign infoMetaMem_tableAid_MPORT_259_data = 6'h0;
  assign infoMetaMem_tableAid_MPORT_259_addr = match_Id;
  assign infoMetaMem_tableAid_MPORT_259_mask = 1'h1;
  assign infoMetaMem_tableAid_MPORT_259_en = _T & _T_1046;
  assign io_tableA_wdata_ready = state == 3'h0; // @[DFCTableD.scala 32:23]
  assign io_tableA_ldata_ready = state == 3'h0; // @[DFCTableD.scala 32:23]
  assign io_tableA_wresp_valid = _T_1058 ? 1'h0 : _GEN_43; // @[Conditional.scala 40:58 DFCTableD.scala 47:25]
  assign io_tableA_wresp_bits = _T_1058 ? 1'h0 : _GEN_44; // @[Conditional.scala 40:58 DFCTableD.scala 48:25]
  assign io_tableA_lresp_valid = _T_1058 ? 1'h0 : _GEN_45; // @[Conditional.scala 40:58 DFCTableD.scala 50:25]
  assign io_tableA_lresp_bits_tableAId = cDown_Id == 6'h0 ? cDown_Id_reg : cDown_Id; // @[DFCTableD.scala 52:39]
  assign io_tableA_lresp_bits_finish = _T_1058 | _GEN_46; // @[Conditional.scala 40:58 DFCTableD.scala 51:31]
  always @(posedge clock) begin
    if(addrMetaMem_listenAddr_MPORT_256_en & addrMetaMem_listenAddr_MPORT_256_mask) begin
      addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_256_addr] <= addrMetaMem_listenAddr_MPORT_256_data; // @[DFCTableD.scala 25:32]
    end
    if(addrMetaMem_listenAddr_MPORT_258_en & addrMetaMem_listenAddr_MPORT_258_mask) begin
      addrMetaMem_listenAddr[addrMetaMem_listenAddr_MPORT_258_addr] <= addrMetaMem_listenAddr_MPORT_258_data; // @[DFCTableD.scala 25:32]
    end
    if(infoMetaMem_tableAid_MPORT_257_en & infoMetaMem_tableAid_MPORT_257_mask) begin
      infoMetaMem_tableAid[infoMetaMem_tableAid_MPORT_257_addr] <= infoMetaMem_tableAid_MPORT_257_data; // @[DFCTableD.scala 26:32]
    end
    if(infoMetaMem_tableAid_MPORT_259_en & infoMetaMem_tableAid_MPORT_259_mask) begin
      infoMetaMem_tableAid[infoMetaMem_tableAid_MPORT_259_addr] <= infoMetaMem_tableAid_MPORT_259_data; // @[DFCTableD.scala 26:32]
    end
    if (_T_1028) begin
      infoMetaMem_tableAid_MPORT_255_addr_pipe_0 <= 8'hff;
    end else if (laddr_reg == addrMetaMem_listenAddr_MPORT_253_data) begin // @[DFCTableD.scala 72:21]
      infoMetaMem_tableAid_MPORT_255_addr_pipe_0 <= 8'hfe;
    end else if (laddr_reg == addrMetaMem_listenAddr_MPORT_252_data) begin // @[DFCTableD.scala 72:21]
      infoMetaMem_tableAid_MPORT_255_addr_pipe_0 <= 8'hfd;
    end else if (laddr_reg == addrMetaMem_listenAddr_MPORT_251_data) begin // @[DFCTableD.scala 72:21]
      infoMetaMem_tableAid_MPORT_255_addr_pipe_0 <= 8'hfc;
    end else begin
      infoMetaMem_tableAid_MPORT_255_addr_pipe_0 <= _T_1021;
    end
    if (reset) begin // @[DFCTableD.scala 27:29]
      tableD_valid <= 256'h0; // @[DFCTableD.scala 27:29]
    end else if (_T & laststate != 3'h5) begin // @[DFCTableD.scala 96:53]
      tableD_valid <= _T_1052; // @[DFCTableD.scala 99:18]
    end else if (state == 3'h1) begin // @[DFCTableD.scala 89:26]
      tableD_valid <= _T_1036; // @[DFCTableD.scala 92:18]
    end
    if (reset) begin // @[DFCTableD.scala 30:22]
      state <= 3'h0; // @[DFCTableD.scala 30:22]
    end else if (_T_1058) begin // @[Conditional.scala 40:58]
      if (io_tableA_wdata_valid) begin // @[DFCTableD.scala 107:34]
        state <= 3'h1; // @[DFCTableD.scala 108:15]
      end else if (io_tableA_ldata_valid) begin // @[DFCTableD.scala 109:40]
        state <= 3'h3; // @[DFCTableD.scala 110:15]
      end
    end else if (_T_1059) begin // @[Conditional.scala 39:67]
      state <= 3'h2; // @[DFCTableD.scala 114:13]
    end else if (_T_1060) begin // @[Conditional.scala 39:67]
      state <= _GEN_22;
    end else begin
      state <= _GEN_34;
    end
    laststate <= state; // @[DFCTableD.scala 31:26]
    if (reset) begin // @[DFCTableD.scala 35:26]
      laddr_reg <= 32'h0; // @[DFCTableD.scala 35:26]
    end else if (is_idle & io_tableA_ldata_valid) begin // @[DFCTableD.scala 65:41]
      laddr_reg <= io_tableA_ldata_bits_listenAddr; // @[DFCTableD.scala 66:15]
    end else if (is_idle & io_tableA_wdata_valid) begin // @[DFCTableD.scala 60:41]
      laddr_reg <= io_tableA_wdata_bits_listenAddr; // @[DFCTableD.scala 61:15]
    end
    if (reset) begin // @[DFCTableD.scala 36:29]
      tableAid_reg <= 6'h0; // @[DFCTableD.scala 36:29]
    end else if (is_idle & io_tableA_wdata_valid) begin // @[DFCTableD.scala 60:41]
      tableAid_reg <= io_tableA_wdata_bits_tableAId; // @[DFCTableD.scala 62:18]
    end
    if (reset) begin // @[DFCTableD.scala 37:26]
      tableD_Id <= 8'h1; // @[DFCTableD.scala 37:26]
    end else if (is_idle & io_tableA_wdata_valid) begin // @[DFCTableD.scala 60:41]
      if (tableD_valid[255]) begin // @[DFCTableD.scala 57:21]
        if (tableD_valid[254]) begin // @[DFCTableD.scala 57:21]
          tableD_Id <= _T_511;
        end else begin
          tableD_Id <= 8'hfe;
        end
      end else begin
        tableD_Id <= 8'hff;
      end
    end
    if (reset) begin // @[DFCTableD.scala 38:25]
      match_Id <= 8'h1; // @[DFCTableD.scala 38:25]
    end else if (state == 3'h3) begin // @[DFCTableD.scala 74:26]
      if (laddr_reg == addrMetaMem_listenAddr_MPORT_254_data) begin // @[DFCTableD.scala 72:21]
        match_Id <= 8'hff;
      end else if (laddr_reg == addrMetaMem_listenAddr_MPORT_253_data) begin // @[DFCTableD.scala 72:21]
        match_Id <= 8'hfe;
      end else begin
        match_Id <= _T_1025;
      end
    end
    if (reset) begin // @[DFCTableD.scala 39:25]
      cDown_Id <= 6'h1; // @[DFCTableD.scala 39:25]
    end else begin
      cDown_Id <= infoMetaMem_tableAid_MPORT_255_data; // @[DFCTableD.scala 78:12]
    end
    if (reset) begin // @[DFCTableD.scala 40:29]
      cDown_Id_reg <= 6'h1; // @[DFCTableD.scala 40:29]
    end else if (state == 3'h5) begin // @[DFCTableD.scala 41:22]
      if (laststate == 3'h4) begin // @[DFCTableD.scala 41:44]
        cDown_Id_reg <= cDown_Id;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1034 & ~reset) begin
          $fwrite(32'h80000002,"[WTD](id: %d).addrMeta.listenAddr = %x\n",tableD_Id,laddr_reg); // @[DFCTableD.scala 93:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1034 & _T_1042) begin
          $fwrite(32'h80000002,"[WTD](id: %d).infoMeta.tableAid = %d\n",tableD_Id,tableAid_reg); // @[DFCTableD.scala 94:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1042) begin
          $fwrite(32'h80000002,"[LTD](id: %d).addrMeta.listenAddr init\n",match_Id); // @[DFCTableD.scala 100:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1047 & _T_1042) begin
          $fwrite(32'h80000002,"[LTD](id: %d).infoMeta.tableAid init\n",match_Id); // @[DFCTableD.scala 101:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    addrMetaMem_listenAddr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    infoMetaMem_tableAid[initvar] = _RAND_1[5:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  infoMetaMem_tableAid_MPORT_255_addr_pipe_0 = _RAND_2[7:0];
  _RAND_3 = {8{`RANDOM}};
  tableD_valid = _RAND_3[255:0];
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  laststate = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  laddr_reg = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  tableAid_reg = _RAND_7[5:0];
  _RAND_8 = {1{`RANDOM}};
  tableD_Id = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  match_Id = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  cDown_Id = _RAND_10[5:0];
  _RAND_11 = {1{`RANDOM}};
  cDown_Id_reg = _RAND_11[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DFCArbiter(
  output        io_cpu1_w_data_ready,
  input         io_cpu1_w_data_valid,
  input  [31:0] io_cpu1_w_data_bits_listenAddr,
  input  [15:0] io_cpu1_w_data_bits_wPid,
  output        io_cpu2_w_data_ready,
  input         io_cpu2_w_data_valid,
  input  [31:0] io_cpu2_w_data_bits_listenAddr,
  input  [15:0] io_cpu2_w_data_bits_wPid,
  output        io_cpu1_l_data_ready,
  input         io_cpu1_l_data_valid,
  input  [31:0] io_cpu1_l_data_bits_listenAddr,
  output        io_cpu2_l_data_ready,
  input         io_cpu2_l_data_valid,
  input  [31:0] io_cpu2_l_data_bits_listenAddr,
  input         io_table_w_data_ready,
  output        io_table_w_data_valid,
  output [31:0] io_table_w_data_bits_listenAddr,
  output [15:0] io_table_w_data_bits_wPid,
  input         io_table_l_data_ready,
  output        io_table_l_data_valid,
  output [31:0] io_table_l_data_bits_listenAddr
);
  wire  _T_6 = ~io_table_w_data_valid; // @[DFCArbiter.scala 33:78]
  assign io_cpu1_w_data_ready = io_table_w_data_ready; // @[DFCArbiter.scala 23:24]
  assign io_cpu2_w_data_ready = io_cpu1_w_data_ready & ~io_cpu1_w_data_valid; // @[DFCArbiter.scala 24:48]
  assign io_cpu1_l_data_ready = io_table_l_data_ready & _T_6; // @[DFCArbiter.scala 34:49]
  assign io_cpu2_l_data_ready = io_cpu1_l_data_ready & ~io_cpu1_l_data_valid; // @[DFCArbiter.scala 35:48]
  assign io_table_w_data_valid = io_cpu1_w_data_valid | io_cpu2_w_data_valid; // @[DFCArbiter.scala 22:50]
  assign io_table_w_data_bits_listenAddr = io_cpu1_w_data_valid ? io_cpu1_w_data_bits_listenAddr :
    io_cpu2_w_data_bits_listenAddr; // @[DFCArbiter.scala 25:41]
  assign io_table_w_data_bits_wPid = io_cpu1_w_data_valid ? io_cpu1_w_data_bits_wPid : io_cpu2_w_data_bits_wPid; // @[DFCArbiter.scala 28:35]
  assign io_table_l_data_valid = (io_cpu1_l_data_valid | io_cpu2_l_data_valid) & ~io_table_w_data_valid; // @[DFCArbiter.scala 33:75]
  assign io_table_l_data_bits_listenAddr = io_cpu1_l_data_valid ? io_cpu1_l_data_bits_listenAddr :
    io_cpu2_l_data_bits_listenAddr; // @[DFCArbiter.scala 36:41]
endmodule
module MemFifo(
  input         clock,
  input         reset,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_listenAddr,
  input  [15:0] io_enq_bits_wPid,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_listenAddr,
  output [15:0] io_deq_bits_wPid
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem_listenAddr [0:7]; // @[DFCfifo.scala 28:25]
  wire [31:0] mem_listenAddr_data_data; // @[DFCfifo.scala 28:25]
  wire [2:0] mem_listenAddr_data_addr; // @[DFCfifo.scala 28:25]
  wire [31:0] mem_listenAddr_MPORT_data; // @[DFCfifo.scala 28:25]
  wire [2:0] mem_listenAddr_MPORT_addr; // @[DFCfifo.scala 28:25]
  wire  mem_listenAddr_MPORT_mask; // @[DFCfifo.scala 28:25]
  wire  mem_listenAddr_MPORT_en; // @[DFCfifo.scala 28:25]
  reg  mem_listenAddr_data_en_pipe_0;
  reg [2:0] mem_listenAddr_data_addr_pipe_0;
  reg [15:0] mem_wPid [0:7]; // @[DFCfifo.scala 28:25]
  wire [15:0] mem_wPid_data_data; // @[DFCfifo.scala 28:25]
  wire [2:0] mem_wPid_data_addr; // @[DFCfifo.scala 28:25]
  wire [15:0] mem_wPid_MPORT_data; // @[DFCfifo.scala 28:25]
  wire [2:0] mem_wPid_MPORT_addr; // @[DFCfifo.scala 28:25]
  wire  mem_wPid_MPORT_mask; // @[DFCfifo.scala 28:25]
  wire  mem_wPid_MPORT_en; // @[DFCfifo.scala 28:25]
  reg  mem_wPid_data_en_pipe_0;
  reg [2:0] mem_wPid_data_addr_pipe_0;
  reg [2:0] readPtr; // @[DFCfifo.scala 20:26]
  wire [2:0] _T_2 = readPtr + 3'h1; // @[DFCfifo.scala 21:60]
  wire [2:0] nextRead = readPtr == 3'h7 ? 3'h0 : _T_2; // @[DFCfifo.scala 21:22]
  reg [1:0] stateReg; // @[DFCfifo.scala 39:25]
  wire  _T_9 = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  reg  emptyReg; // @[DFCfifo.scala 35:25]
  wire  _T_10 = ~emptyReg; // @[DFCfifo.scala 55:13]
  wire  _T_12 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _GEN_22 = io_deq_ready & _T_10; // @[DFCfifo.scala 63:26]
  wire  _T_15 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _GEN_40 = _T_12 ? _GEN_22 : _T_15 & _GEN_22; // @[Conditional.scala 39:67]
  wire  incrRead = _T_9 ? _T_10 : _GEN_40; // @[Conditional.scala 40:58]
  reg [2:0] writePtr; // @[DFCfifo.scala 20:26]
  wire [2:0] _T_5 = writePtr + 3'h1; // @[DFCfifo.scala 21:60]
  wire [2:0] nextWrite = writePtr == 3'h7 ? 3'h0 : _T_5; // @[DFCfifo.scala 21:22]
  reg  fullReg; // @[DFCfifo.scala 36:24]
  wire  _T_6 = ~fullReg; // @[DFCfifo.scala 42:25]
  wire  incrWrite = io_enq_valid & ~fullReg; // @[DFCfifo.scala 42:22]
  reg [31:0] shadowReg_listenAddr; // @[DFCfifo.scala 41:22]
  reg [15:0] shadowReg_wPid; // @[DFCfifo.scala 41:22]
  wire  _GEN_9 = incrWrite ? 1'h0 : emptyReg; // @[DFCfifo.scala 42:35 DFCfifo.scala 44:14 DFCfifo.scala 35:25]
  wire  _GEN_10 = incrWrite ? nextWrite == readPtr : fullReg; // @[DFCfifo.scala 42:35 DFCfifo.scala 45:13 DFCfifo.scala 36:24]
  wire  _GEN_12 = ~emptyReg ? 1'h0 : _GEN_10; // @[DFCfifo.scala 55:24 DFCfifo.scala 57:17]
  wire  _GEN_13 = ~emptyReg ? nextRead == writePtr : _GEN_9; // @[DFCfifo.scala 55:24 DFCfifo.scala 58:18]
  wire [1:0] _GEN_15 = _T_10 ? 2'h1 : 2'h0; // @[DFCfifo.scala 64:27 DFCfifo.scala 65:20 DFCfifo.scala 70:20]
  wire  _GEN_20 = io_deq_ready ? _GEN_12 : _GEN_10; // @[DFCfifo.scala 63:26]
  wire  _GEN_21 = io_deq_ready ? _GEN_13 : _GEN_9; // @[DFCfifo.scala 63:26]
  wire [1:0] _GEN_29 = io_deq_ready ? _GEN_15 : stateReg; // @[DFCfifo.scala 78:26 DFCfifo.scala 39:25]
  wire  _GEN_35 = _T_15 ? _GEN_21 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_39 = _T_12 ? _GEN_21 : _GEN_35; // @[Conditional.scala 39:67]
  wire  _GEN_45 = _T_9 ? _GEN_13 : _GEN_39; // @[Conditional.scala 40:58]
  wire  _T_18 = stateReg == 2'h1; // @[DFCfifo.scala 90:31]
  assign mem_listenAddr_data_addr = mem_listenAddr_data_addr_pipe_0;
  assign mem_listenAddr_data_data = mem_listenAddr[mem_listenAddr_data_addr]; // @[DFCfifo.scala 28:25]
  assign mem_listenAddr_MPORT_data = io_enq_bits_listenAddr;
  assign mem_listenAddr_MPORT_addr = writePtr;
  assign mem_listenAddr_MPORT_mask = 1'h1;
  assign mem_listenAddr_MPORT_en = io_enq_valid & _T_6;
  assign mem_wPid_data_addr = mem_wPid_data_addr_pipe_0;
  assign mem_wPid_data_data = mem_wPid[mem_wPid_data_addr]; // @[DFCfifo.scala 28:25]
  assign mem_wPid_MPORT_data = io_enq_bits_wPid;
  assign mem_wPid_MPORT_addr = writePtr;
  assign mem_wPid_MPORT_mask = 1'h1;
  assign mem_wPid_MPORT_en = io_enq_valid & _T_6;
  assign io_deq_valid = _T_18 | stateReg == 2'h2; // @[DFCfifo.scala 92:38]
  assign io_deq_bits_listenAddr = stateReg == 2'h1 ? mem_listenAddr_data_data : shadowReg_listenAddr; // @[DFCfifo.scala 90:21]
  assign io_deq_bits_wPid = stateReg == 2'h1 ? mem_wPid_data_data : shadowReg_wPid; // @[DFCfifo.scala 90:21]
  always @(posedge clock) begin
    if(mem_listenAddr_MPORT_en & mem_listenAddr_MPORT_mask) begin
      mem_listenAddr[mem_listenAddr_MPORT_addr] <= mem_listenAddr_MPORT_data; // @[DFCfifo.scala 28:25]
    end
    if (_T_9) begin
      mem_listenAddr_data_en_pipe_0 <= _T_10;
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      mem_listenAddr_data_en_pipe_0 <= _GEN_22;
    end else begin
      mem_listenAddr_data_en_pipe_0 <= _T_15 & _GEN_22;
    end
    if (_T_9 ? _T_10 : _GEN_40) begin
      mem_listenAddr_data_addr_pipe_0 <= readPtr;
    end
    if(mem_wPid_MPORT_en & mem_wPid_MPORT_mask) begin
      mem_wPid[mem_wPid_MPORT_addr] <= mem_wPid_MPORT_data; // @[DFCfifo.scala 28:25]
    end
    if (_T_9) begin
      mem_wPid_data_en_pipe_0 <= _T_10;
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      mem_wPid_data_en_pipe_0 <= _GEN_22;
    end else begin
      mem_wPid_data_en_pipe_0 <= _T_15 & _GEN_22;
    end
    if (_T_9 ? _T_10 : _GEN_40) begin
      mem_wPid_data_addr_pipe_0 <= readPtr;
    end
    if (reset) begin // @[DFCfifo.scala 20:26]
      readPtr <= 3'h0; // @[DFCfifo.scala 20:26]
    end else if (incrRead) begin // @[DFCfifo.scala 22:17]
      if (readPtr == 3'h7) begin // @[DFCfifo.scala 21:22]
        readPtr <= 3'h0;
      end else begin
        readPtr <= _T_2;
      end
    end
    if (reset) begin // @[DFCfifo.scala 39:25]
      stateReg <= 2'h0; // @[DFCfifo.scala 39:25]
    end else if (_T_9) begin // @[Conditional.scala 40:58]
      if (~emptyReg) begin // @[DFCfifo.scala 55:24]
        stateReg <= 2'h1; // @[DFCfifo.scala 56:18]
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (io_deq_ready) begin // @[DFCfifo.scala 63:26]
        stateReg <= _GEN_15;
      end else begin
        stateReg <= 2'h2; // @[DFCfifo.scala 74:18]
      end
    end else if (_T_15) begin // @[Conditional.scala 39:67]
      stateReg <= _GEN_29;
    end
    emptyReg <= reset | _GEN_45; // @[DFCfifo.scala 35:25 DFCfifo.scala 35:25]
    if (reset) begin // @[DFCfifo.scala 20:26]
      writePtr <= 3'h0; // @[DFCfifo.scala 20:26]
    end else if (incrWrite) begin // @[DFCfifo.scala 22:17]
      if (writePtr == 3'h7) begin // @[DFCfifo.scala 21:22]
        writePtr <= 3'h0;
      end else begin
        writePtr <= _T_5;
      end
    end
    if (reset) begin // @[DFCfifo.scala 36:24]
      fullReg <= 1'h0; // @[DFCfifo.scala 36:24]
    end else if (_T_9) begin // @[Conditional.scala 40:58]
      fullReg <= _GEN_12;
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      fullReg <= _GEN_20;
    end else if (_T_15) begin // @[Conditional.scala 39:67]
      fullReg <= _GEN_20;
    end else begin
      fullReg <= _GEN_10;
    end
    if (!(_T_9)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (!(io_deq_ready)) begin // @[DFCfifo.scala 63:26]
          shadowReg_listenAddr <= mem_listenAddr_data_data; // @[DFCfifo.scala 73:19]
        end
      end
    end
    if (!(_T_9)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (!(io_deq_ready)) begin // @[DFCfifo.scala 63:26]
          shadowReg_wPid <= mem_wPid_data_data; // @[DFCfifo.scala 73:19]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    mem_listenAddr[initvar] = _RAND_0[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    mem_wPid[initvar] = _RAND_3[15:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_listenAddr_data_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_listenAddr_data_addr_pipe_0 = _RAND_2[2:0];
  _RAND_4 = {1{`RANDOM}};
  mem_wPid_data_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  mem_wPid_data_addr_pipe_0 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  readPtr = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  stateReg = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  emptyReg = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  writePtr = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  fullReg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  shadowReg_listenAddr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  shadowReg_wPid = _RAND_12[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemFifo_2(
  input         clock,
  input         reset,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_listenAddr,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_listenAddr
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mem_listenAddr [0:7]; // @[DFCfifo.scala 28:25]
  wire [31:0] mem_listenAddr_data_data; // @[DFCfifo.scala 28:25]
  wire [2:0] mem_listenAddr_data_addr; // @[DFCfifo.scala 28:25]
  wire [31:0] mem_listenAddr_MPORT_data; // @[DFCfifo.scala 28:25]
  wire [2:0] mem_listenAddr_MPORT_addr; // @[DFCfifo.scala 28:25]
  wire  mem_listenAddr_MPORT_mask; // @[DFCfifo.scala 28:25]
  wire  mem_listenAddr_MPORT_en; // @[DFCfifo.scala 28:25]
  reg  mem_listenAddr_data_en_pipe_0;
  reg [2:0] mem_listenAddr_data_addr_pipe_0;
  reg [2:0] readPtr; // @[DFCfifo.scala 20:26]
  wire [2:0] _T_2 = readPtr + 3'h1; // @[DFCfifo.scala 21:60]
  wire [2:0] nextRead = readPtr == 3'h7 ? 3'h0 : _T_2; // @[DFCfifo.scala 21:22]
  reg [1:0] stateReg; // @[DFCfifo.scala 39:25]
  wire  _T_9 = 2'h0 == stateReg; // @[Conditional.scala 37:30]
  reg  emptyReg; // @[DFCfifo.scala 35:25]
  wire  _T_10 = ~emptyReg; // @[DFCfifo.scala 55:13]
  wire  _T_12 = 2'h1 == stateReg; // @[Conditional.scala 37:30]
  wire  _GEN_21 = io_deq_ready & _T_10; // @[DFCfifo.scala 63:26]
  wire  _T_15 = 2'h2 == stateReg; // @[Conditional.scala 37:30]
  wire  _GEN_38 = _T_12 ? _GEN_21 : _T_15 & _GEN_21; // @[Conditional.scala 39:67]
  wire  incrRead = _T_9 ? _T_10 : _GEN_38; // @[Conditional.scala 40:58]
  reg [2:0] writePtr; // @[DFCfifo.scala 20:26]
  wire [2:0] _T_5 = writePtr + 3'h1; // @[DFCfifo.scala 21:60]
  wire [2:0] nextWrite = writePtr == 3'h7 ? 3'h0 : _T_5; // @[DFCfifo.scala 21:22]
  reg  fullReg; // @[DFCfifo.scala 36:24]
  wire  _T_6 = ~fullReg; // @[DFCfifo.scala 42:25]
  wire  incrWrite = io_enq_valid & ~fullReg; // @[DFCfifo.scala 42:22]
  reg [31:0] shadowReg_listenAddr; // @[DFCfifo.scala 41:22]
  wire  _GEN_8 = incrWrite ? 1'h0 : emptyReg; // @[DFCfifo.scala 42:35 DFCfifo.scala 44:14 DFCfifo.scala 35:25]
  wire  _GEN_9 = incrWrite ? nextWrite == readPtr : fullReg; // @[DFCfifo.scala 42:35 DFCfifo.scala 45:13 DFCfifo.scala 36:24]
  wire  _GEN_11 = ~emptyReg ? 1'h0 : _GEN_9; // @[DFCfifo.scala 55:24 DFCfifo.scala 57:17]
  wire  _GEN_12 = ~emptyReg ? nextRead == writePtr : _GEN_8; // @[DFCfifo.scala 55:24 DFCfifo.scala 58:18]
  wire [1:0] _GEN_14 = _T_10 ? 2'h1 : 2'h0; // @[DFCfifo.scala 64:27 DFCfifo.scala 65:20 DFCfifo.scala 70:20]
  wire  _GEN_19 = io_deq_ready ? _GEN_11 : _GEN_9; // @[DFCfifo.scala 63:26]
  wire  _GEN_20 = io_deq_ready ? _GEN_12 : _GEN_8; // @[DFCfifo.scala 63:26]
  wire [1:0] _GEN_27 = io_deq_ready ? _GEN_14 : stateReg; // @[DFCfifo.scala 78:26 DFCfifo.scala 39:25]
  wire  _GEN_33 = _T_15 ? _GEN_20 : _GEN_8; // @[Conditional.scala 39:67]
  wire  _GEN_37 = _T_12 ? _GEN_20 : _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_9 ? _GEN_12 : _GEN_37; // @[Conditional.scala 40:58]
  wire  _T_18 = stateReg == 2'h1; // @[DFCfifo.scala 90:31]
  assign mem_listenAddr_data_addr = mem_listenAddr_data_addr_pipe_0;
  assign mem_listenAddr_data_data = mem_listenAddr[mem_listenAddr_data_addr]; // @[DFCfifo.scala 28:25]
  assign mem_listenAddr_MPORT_data = io_enq_bits_listenAddr;
  assign mem_listenAddr_MPORT_addr = writePtr;
  assign mem_listenAddr_MPORT_mask = 1'h1;
  assign mem_listenAddr_MPORT_en = io_enq_valid & _T_6;
  assign io_deq_valid = _T_18 | stateReg == 2'h2; // @[DFCfifo.scala 92:38]
  assign io_deq_bits_listenAddr = stateReg == 2'h1 ? mem_listenAddr_data_data : shadowReg_listenAddr; // @[DFCfifo.scala 90:21]
  always @(posedge clock) begin
    if(mem_listenAddr_MPORT_en & mem_listenAddr_MPORT_mask) begin
      mem_listenAddr[mem_listenAddr_MPORT_addr] <= mem_listenAddr_MPORT_data; // @[DFCfifo.scala 28:25]
    end
    if (_T_9) begin
      mem_listenAddr_data_en_pipe_0 <= _T_10;
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      mem_listenAddr_data_en_pipe_0 <= _GEN_21;
    end else begin
      mem_listenAddr_data_en_pipe_0 <= _T_15 & _GEN_21;
    end
    if (_T_9 ? _T_10 : _GEN_38) begin
      mem_listenAddr_data_addr_pipe_0 <= readPtr;
    end
    if (reset) begin // @[DFCfifo.scala 20:26]
      readPtr <= 3'h0; // @[DFCfifo.scala 20:26]
    end else if (incrRead) begin // @[DFCfifo.scala 22:17]
      if (readPtr == 3'h7) begin // @[DFCfifo.scala 21:22]
        readPtr <= 3'h0;
      end else begin
        readPtr <= _T_2;
      end
    end
    if (reset) begin // @[DFCfifo.scala 39:25]
      stateReg <= 2'h0; // @[DFCfifo.scala 39:25]
    end else if (_T_9) begin // @[Conditional.scala 40:58]
      if (~emptyReg) begin // @[DFCfifo.scala 55:24]
        stateReg <= 2'h1; // @[DFCfifo.scala 56:18]
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      if (io_deq_ready) begin // @[DFCfifo.scala 63:26]
        stateReg <= _GEN_14;
      end else begin
        stateReg <= 2'h2; // @[DFCfifo.scala 74:18]
      end
    end else if (_T_15) begin // @[Conditional.scala 39:67]
      stateReg <= _GEN_27;
    end
    emptyReg <= reset | _GEN_42; // @[DFCfifo.scala 35:25 DFCfifo.scala 35:25]
    if (reset) begin // @[DFCfifo.scala 20:26]
      writePtr <= 3'h0; // @[DFCfifo.scala 20:26]
    end else if (incrWrite) begin // @[DFCfifo.scala 22:17]
      if (writePtr == 3'h7) begin // @[DFCfifo.scala 21:22]
        writePtr <= 3'h0;
      end else begin
        writePtr <= _T_5;
      end
    end
    if (reset) begin // @[DFCfifo.scala 36:24]
      fullReg <= 1'h0; // @[DFCfifo.scala 36:24]
    end else if (_T_9) begin // @[Conditional.scala 40:58]
      fullReg <= _GEN_11;
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      fullReg <= _GEN_19;
    end else if (_T_15) begin // @[Conditional.scala 39:67]
      fullReg <= _GEN_19;
    end else begin
      fullReg <= _GEN_9;
    end
    if (!(_T_9)) begin // @[Conditional.scala 40:58]
      if (_T_12) begin // @[Conditional.scala 39:67]
        if (!(io_deq_ready)) begin // @[DFCfifo.scala 63:26]
          shadowReg_listenAddr <= mem_listenAddr_data_data; // @[DFCfifo.scala 73:19]
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    mem_listenAddr[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_listenAddr_data_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_listenAddr_data_addr_pipe_0 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  readPtr = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  stateReg = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  emptyReg = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  writePtr = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  fullReg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  shadowReg_listenAddr = _RAND_8[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DFCExptArbiter(
  output        io_table_e_data_ready,
  input         io_table_e_data_valid,
  input  [15:0] io_table_e_data_bits_pid,
  input         io_cpu1_e_data_ready,
  output        io_cpu1_e_data_valid,
  output [15:0] io_cpu1_e_data_bits_pid
);
  assign io_table_e_data_ready = io_cpu1_e_data_ready; // @[DFCTable.scala 97:49]
  assign io_cpu1_e_data_valid = io_table_e_data_valid & io_cpu1_e_data_ready; // @[DFCTable.scala 98:49]
  assign io_cpu1_e_data_bits_pid = io_table_e_data_bits_pid; // @[DFCTable.scala 95:23]
endmodule
module DFC_Table(
  input         clock,
  input         reset,
  input         io_cpu1_w_data_valid,
  input  [31:0] io_cpu1_w_data_bits_listenAddr,
  input  [15:0] io_cpu1_w_data_bits_wPid,
  input         io_cpu1_l_data_valid,
  input  [31:0] io_cpu1_l_data_bits_listenAddr,
  input         io_cpu1_e_data_ready,
  output        io_cpu1_e_data_valid,
  output [15:0] io_cpu1_e_data_bits_pid,
  output        io_cpu_f_data_valid,
  output        io_cpu_f_data_bits_full_sig
);
  wire  dfc_tableA_clock; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_reset; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_cpu_w_data_ready; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_cpu_w_data_valid; // @[DFCTable.scala 108:26]
  wire [31:0] dfc_tableA_io_cpu_w_data_bits_listenAddr; // @[DFCTable.scala 108:26]
  wire [15:0] dfc_tableA_io_cpu_w_data_bits_wPid; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_cpu_l_data_ready; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_cpu_l_data_valid; // @[DFCTable.scala 108:26]
  wire [31:0] dfc_tableA_io_cpu_l_data_bits_listenAddr; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_tableD_wdata_ready; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_tableD_wdata_valid; // @[DFCTable.scala 108:26]
  wire [31:0] dfc_tableA_io_tableD_wdata_bits_listenAddr; // @[DFCTable.scala 108:26]
  wire [5:0] dfc_tableA_io_tableD_wdata_bits_tableAId; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_tableD_ldata_ready; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_tableD_ldata_valid; // @[DFCTable.scala 108:26]
  wire [31:0] dfc_tableA_io_tableD_ldata_bits_listenAddr; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_tableD_wresp_ready; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_tableD_wresp_valid; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_tableD_wresp_bits; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_tableD_lresp_ready; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_tableD_lresp_valid; // @[DFCTable.scala 108:26]
  wire [5:0] dfc_tableA_io_tableD_lresp_bits_tableAId; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_tableD_lresp_bits_finish; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_cpu_expt_data_ready; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_cpu_expt_data_valid; // @[DFCTable.scala 108:26]
  wire [15:0] dfc_tableA_io_cpu_expt_data_bits_pid; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_dfc_full_data_valid; // @[DFCTable.scala 108:26]
  wire  dfc_tableA_io_dfc_full_data_bits_full_sig; // @[DFCTable.scala 108:26]
  wire  dfc_tableD_clock; // @[DFCTable.scala 109:26]
  wire  dfc_tableD_reset; // @[DFCTable.scala 109:26]
  wire  dfc_tableD_io_tableA_wdata_ready; // @[DFCTable.scala 109:26]
  wire  dfc_tableD_io_tableA_wdata_valid; // @[DFCTable.scala 109:26]
  wire [31:0] dfc_tableD_io_tableA_wdata_bits_listenAddr; // @[DFCTable.scala 109:26]
  wire [5:0] dfc_tableD_io_tableA_wdata_bits_tableAId; // @[DFCTable.scala 109:26]
  wire  dfc_tableD_io_tableA_ldata_ready; // @[DFCTable.scala 109:26]
  wire  dfc_tableD_io_tableA_ldata_valid; // @[DFCTable.scala 109:26]
  wire [31:0] dfc_tableD_io_tableA_ldata_bits_listenAddr; // @[DFCTable.scala 109:26]
  wire  dfc_tableD_io_tableA_wresp_ready; // @[DFCTable.scala 109:26]
  wire  dfc_tableD_io_tableA_wresp_valid; // @[DFCTable.scala 109:26]
  wire  dfc_tableD_io_tableA_wresp_bits; // @[DFCTable.scala 109:26]
  wire  dfc_tableD_io_tableA_lresp_ready; // @[DFCTable.scala 109:26]
  wire  dfc_tableD_io_tableA_lresp_valid; // @[DFCTable.scala 109:26]
  wire [5:0] dfc_tableD_io_tableA_lresp_bits_tableAId; // @[DFCTable.scala 109:26]
  wire  dfc_tableD_io_tableA_lresp_bits_finish; // @[DFCTable.scala 109:26]
  wire  dfc_arbiter_io_cpu1_w_data_ready; // @[DFCTable.scala 110:27]
  wire  dfc_arbiter_io_cpu1_w_data_valid; // @[DFCTable.scala 110:27]
  wire [31:0] dfc_arbiter_io_cpu1_w_data_bits_listenAddr; // @[DFCTable.scala 110:27]
  wire [15:0] dfc_arbiter_io_cpu1_w_data_bits_wPid; // @[DFCTable.scala 110:27]
  wire  dfc_arbiter_io_cpu2_w_data_ready; // @[DFCTable.scala 110:27]
  wire  dfc_arbiter_io_cpu2_w_data_valid; // @[DFCTable.scala 110:27]
  wire [31:0] dfc_arbiter_io_cpu2_w_data_bits_listenAddr; // @[DFCTable.scala 110:27]
  wire [15:0] dfc_arbiter_io_cpu2_w_data_bits_wPid; // @[DFCTable.scala 110:27]
  wire  dfc_arbiter_io_cpu1_l_data_ready; // @[DFCTable.scala 110:27]
  wire  dfc_arbiter_io_cpu1_l_data_valid; // @[DFCTable.scala 110:27]
  wire [31:0] dfc_arbiter_io_cpu1_l_data_bits_listenAddr; // @[DFCTable.scala 110:27]
  wire  dfc_arbiter_io_cpu2_l_data_ready; // @[DFCTable.scala 110:27]
  wire  dfc_arbiter_io_cpu2_l_data_valid; // @[DFCTable.scala 110:27]
  wire [31:0] dfc_arbiter_io_cpu2_l_data_bits_listenAddr; // @[DFCTable.scala 110:27]
  wire  dfc_arbiter_io_table_w_data_ready; // @[DFCTable.scala 110:27]
  wire  dfc_arbiter_io_table_w_data_valid; // @[DFCTable.scala 110:27]
  wire [31:0] dfc_arbiter_io_table_w_data_bits_listenAddr; // @[DFCTable.scala 110:27]
  wire [15:0] dfc_arbiter_io_table_w_data_bits_wPid; // @[DFCTable.scala 110:27]
  wire  dfc_arbiter_io_table_l_data_ready; // @[DFCTable.scala 110:27]
  wire  dfc_arbiter_io_table_l_data_valid; // @[DFCTable.scala 110:27]
  wire [31:0] dfc_arbiter_io_table_l_data_bits_listenAddr; // @[DFCTable.scala 110:27]
  wire  cpu1_wbuf_clock; // @[DFCTable.scala 111:25]
  wire  cpu1_wbuf_reset; // @[DFCTable.scala 111:25]
  wire  cpu1_wbuf_io_enq_valid; // @[DFCTable.scala 111:25]
  wire [31:0] cpu1_wbuf_io_enq_bits_listenAddr; // @[DFCTable.scala 111:25]
  wire [15:0] cpu1_wbuf_io_enq_bits_wPid; // @[DFCTable.scala 111:25]
  wire  cpu1_wbuf_io_deq_ready; // @[DFCTable.scala 111:25]
  wire  cpu1_wbuf_io_deq_valid; // @[DFCTable.scala 111:25]
  wire [31:0] cpu1_wbuf_io_deq_bits_listenAddr; // @[DFCTable.scala 111:25]
  wire [15:0] cpu1_wbuf_io_deq_bits_wPid; // @[DFCTable.scala 111:25]
  wire  cpu2_wbuf_clock; // @[DFCTable.scala 112:25]
  wire  cpu2_wbuf_reset; // @[DFCTable.scala 112:25]
  wire  cpu2_wbuf_io_enq_valid; // @[DFCTable.scala 112:25]
  wire [31:0] cpu2_wbuf_io_enq_bits_listenAddr; // @[DFCTable.scala 112:25]
  wire [15:0] cpu2_wbuf_io_enq_bits_wPid; // @[DFCTable.scala 112:25]
  wire  cpu2_wbuf_io_deq_ready; // @[DFCTable.scala 112:25]
  wire  cpu2_wbuf_io_deq_valid; // @[DFCTable.scala 112:25]
  wire [31:0] cpu2_wbuf_io_deq_bits_listenAddr; // @[DFCTable.scala 112:25]
  wire [15:0] cpu2_wbuf_io_deq_bits_wPid; // @[DFCTable.scala 112:25]
  wire  cpu1_lbuf_clock; // @[DFCTable.scala 113:25]
  wire  cpu1_lbuf_reset; // @[DFCTable.scala 113:25]
  wire  cpu1_lbuf_io_enq_valid; // @[DFCTable.scala 113:25]
  wire [31:0] cpu1_lbuf_io_enq_bits_listenAddr; // @[DFCTable.scala 113:25]
  wire  cpu1_lbuf_io_deq_ready; // @[DFCTable.scala 113:25]
  wire  cpu1_lbuf_io_deq_valid; // @[DFCTable.scala 113:25]
  wire [31:0] cpu1_lbuf_io_deq_bits_listenAddr; // @[DFCTable.scala 113:25]
  wire  cpu2_lbuf_clock; // @[DFCTable.scala 114:25]
  wire  cpu2_lbuf_reset; // @[DFCTable.scala 114:25]
  wire  cpu2_lbuf_io_enq_valid; // @[DFCTable.scala 114:25]
  wire [31:0] cpu2_lbuf_io_enq_bits_listenAddr; // @[DFCTable.scala 114:25]
  wire  cpu2_lbuf_io_deq_ready; // @[DFCTable.scala 114:25]
  wire  cpu2_lbuf_io_deq_valid; // @[DFCTable.scala 114:25]
  wire [31:0] cpu2_lbuf_io_deq_bits_listenAddr; // @[DFCTable.scala 114:25]
  wire  expt_arbiter_io_table_e_data_ready; // @[DFCTable.scala 115:28]
  wire  expt_arbiter_io_table_e_data_valid; // @[DFCTable.scala 115:28]
  wire [15:0] expt_arbiter_io_table_e_data_bits_pid; // @[DFCTable.scala 115:28]
  wire  expt_arbiter_io_cpu1_e_data_ready; // @[DFCTable.scala 115:28]
  wire  expt_arbiter_io_cpu1_e_data_valid; // @[DFCTable.scala 115:28]
  wire [15:0] expt_arbiter_io_cpu1_e_data_bits_pid; // @[DFCTable.scala 115:28]
  DFC_TableA dfc_tableA ( // @[DFCTable.scala 108:26]
    .clock(dfc_tableA_clock),
    .reset(dfc_tableA_reset),
    .io_cpu_w_data_ready(dfc_tableA_io_cpu_w_data_ready),
    .io_cpu_w_data_valid(dfc_tableA_io_cpu_w_data_valid),
    .io_cpu_w_data_bits_listenAddr(dfc_tableA_io_cpu_w_data_bits_listenAddr),
    .io_cpu_w_data_bits_wPid(dfc_tableA_io_cpu_w_data_bits_wPid),
    .io_cpu_l_data_ready(dfc_tableA_io_cpu_l_data_ready),
    .io_cpu_l_data_valid(dfc_tableA_io_cpu_l_data_valid),
    .io_cpu_l_data_bits_listenAddr(dfc_tableA_io_cpu_l_data_bits_listenAddr),
    .io_tableD_wdata_ready(dfc_tableA_io_tableD_wdata_ready),
    .io_tableD_wdata_valid(dfc_tableA_io_tableD_wdata_valid),
    .io_tableD_wdata_bits_listenAddr(dfc_tableA_io_tableD_wdata_bits_listenAddr),
    .io_tableD_wdata_bits_tableAId(dfc_tableA_io_tableD_wdata_bits_tableAId),
    .io_tableD_ldata_ready(dfc_tableA_io_tableD_ldata_ready),
    .io_tableD_ldata_valid(dfc_tableA_io_tableD_ldata_valid),
    .io_tableD_ldata_bits_listenAddr(dfc_tableA_io_tableD_ldata_bits_listenAddr),
    .io_tableD_wresp_ready(dfc_tableA_io_tableD_wresp_ready),
    .io_tableD_wresp_valid(dfc_tableA_io_tableD_wresp_valid),
    .io_tableD_wresp_bits(dfc_tableA_io_tableD_wresp_bits),
    .io_tableD_lresp_ready(dfc_tableA_io_tableD_lresp_ready),
    .io_tableD_lresp_valid(dfc_tableA_io_tableD_lresp_valid),
    .io_tableD_lresp_bits_tableAId(dfc_tableA_io_tableD_lresp_bits_tableAId),
    .io_tableD_lresp_bits_finish(dfc_tableA_io_tableD_lresp_bits_finish),
    .io_cpu_expt_data_ready(dfc_tableA_io_cpu_expt_data_ready),
    .io_cpu_expt_data_valid(dfc_tableA_io_cpu_expt_data_valid),
    .io_cpu_expt_data_bits_pid(dfc_tableA_io_cpu_expt_data_bits_pid),
    .io_dfc_full_data_valid(dfc_tableA_io_dfc_full_data_valid),
    .io_dfc_full_data_bits_full_sig(dfc_tableA_io_dfc_full_data_bits_full_sig)
  );
  DFC_TableD dfc_tableD ( // @[DFCTable.scala 109:26]
    .clock(dfc_tableD_clock),
    .reset(dfc_tableD_reset),
    .io_tableA_wdata_ready(dfc_tableD_io_tableA_wdata_ready),
    .io_tableA_wdata_valid(dfc_tableD_io_tableA_wdata_valid),
    .io_tableA_wdata_bits_listenAddr(dfc_tableD_io_tableA_wdata_bits_listenAddr),
    .io_tableA_wdata_bits_tableAId(dfc_tableD_io_tableA_wdata_bits_tableAId),
    .io_tableA_ldata_ready(dfc_tableD_io_tableA_ldata_ready),
    .io_tableA_ldata_valid(dfc_tableD_io_tableA_ldata_valid),
    .io_tableA_ldata_bits_listenAddr(dfc_tableD_io_tableA_ldata_bits_listenAddr),
    .io_tableA_wresp_ready(dfc_tableD_io_tableA_wresp_ready),
    .io_tableA_wresp_valid(dfc_tableD_io_tableA_wresp_valid),
    .io_tableA_wresp_bits(dfc_tableD_io_tableA_wresp_bits),
    .io_tableA_lresp_ready(dfc_tableD_io_tableA_lresp_ready),
    .io_tableA_lresp_valid(dfc_tableD_io_tableA_lresp_valid),
    .io_tableA_lresp_bits_tableAId(dfc_tableD_io_tableA_lresp_bits_tableAId),
    .io_tableA_lresp_bits_finish(dfc_tableD_io_tableA_lresp_bits_finish)
  );
  DFCArbiter dfc_arbiter ( // @[DFCTable.scala 110:27]
    .io_cpu1_w_data_ready(dfc_arbiter_io_cpu1_w_data_ready),
    .io_cpu1_w_data_valid(dfc_arbiter_io_cpu1_w_data_valid),
    .io_cpu1_w_data_bits_listenAddr(dfc_arbiter_io_cpu1_w_data_bits_listenAddr),
    .io_cpu1_w_data_bits_wPid(dfc_arbiter_io_cpu1_w_data_bits_wPid),
    .io_cpu2_w_data_ready(dfc_arbiter_io_cpu2_w_data_ready),
    .io_cpu2_w_data_valid(dfc_arbiter_io_cpu2_w_data_valid),
    .io_cpu2_w_data_bits_listenAddr(dfc_arbiter_io_cpu2_w_data_bits_listenAddr),
    .io_cpu2_w_data_bits_wPid(dfc_arbiter_io_cpu2_w_data_bits_wPid),
    .io_cpu1_l_data_ready(dfc_arbiter_io_cpu1_l_data_ready),
    .io_cpu1_l_data_valid(dfc_arbiter_io_cpu1_l_data_valid),
    .io_cpu1_l_data_bits_listenAddr(dfc_arbiter_io_cpu1_l_data_bits_listenAddr),
    .io_cpu2_l_data_ready(dfc_arbiter_io_cpu2_l_data_ready),
    .io_cpu2_l_data_valid(dfc_arbiter_io_cpu2_l_data_valid),
    .io_cpu2_l_data_bits_listenAddr(dfc_arbiter_io_cpu2_l_data_bits_listenAddr),
    .io_table_w_data_ready(dfc_arbiter_io_table_w_data_ready),
    .io_table_w_data_valid(dfc_arbiter_io_table_w_data_valid),
    .io_table_w_data_bits_listenAddr(dfc_arbiter_io_table_w_data_bits_listenAddr),
    .io_table_w_data_bits_wPid(dfc_arbiter_io_table_w_data_bits_wPid),
    .io_table_l_data_ready(dfc_arbiter_io_table_l_data_ready),
    .io_table_l_data_valid(dfc_arbiter_io_table_l_data_valid),
    .io_table_l_data_bits_listenAddr(dfc_arbiter_io_table_l_data_bits_listenAddr)
  );
  MemFifo cpu1_wbuf ( // @[DFCTable.scala 111:25]
    .clock(cpu1_wbuf_clock),
    .reset(cpu1_wbuf_reset),
    .io_enq_valid(cpu1_wbuf_io_enq_valid),
    .io_enq_bits_listenAddr(cpu1_wbuf_io_enq_bits_listenAddr),
    .io_enq_bits_wPid(cpu1_wbuf_io_enq_bits_wPid),
    .io_deq_ready(cpu1_wbuf_io_deq_ready),
    .io_deq_valid(cpu1_wbuf_io_deq_valid),
    .io_deq_bits_listenAddr(cpu1_wbuf_io_deq_bits_listenAddr),
    .io_deq_bits_wPid(cpu1_wbuf_io_deq_bits_wPid)
  );
  MemFifo cpu2_wbuf ( // @[DFCTable.scala 112:25]
    .clock(cpu2_wbuf_clock),
    .reset(cpu2_wbuf_reset),
    .io_enq_valid(cpu2_wbuf_io_enq_valid),
    .io_enq_bits_listenAddr(cpu2_wbuf_io_enq_bits_listenAddr),
    .io_enq_bits_wPid(cpu2_wbuf_io_enq_bits_wPid),
    .io_deq_ready(cpu2_wbuf_io_deq_ready),
    .io_deq_valid(cpu2_wbuf_io_deq_valid),
    .io_deq_bits_listenAddr(cpu2_wbuf_io_deq_bits_listenAddr),
    .io_deq_bits_wPid(cpu2_wbuf_io_deq_bits_wPid)
  );
  MemFifo_2 cpu1_lbuf ( // @[DFCTable.scala 113:25]
    .clock(cpu1_lbuf_clock),
    .reset(cpu1_lbuf_reset),
    .io_enq_valid(cpu1_lbuf_io_enq_valid),
    .io_enq_bits_listenAddr(cpu1_lbuf_io_enq_bits_listenAddr),
    .io_deq_ready(cpu1_lbuf_io_deq_ready),
    .io_deq_valid(cpu1_lbuf_io_deq_valid),
    .io_deq_bits_listenAddr(cpu1_lbuf_io_deq_bits_listenAddr)
  );
  MemFifo_2 cpu2_lbuf ( // @[DFCTable.scala 114:25]
    .clock(cpu2_lbuf_clock),
    .reset(cpu2_lbuf_reset),
    .io_enq_valid(cpu2_lbuf_io_enq_valid),
    .io_enq_bits_listenAddr(cpu2_lbuf_io_enq_bits_listenAddr),
    .io_deq_ready(cpu2_lbuf_io_deq_ready),
    .io_deq_valid(cpu2_lbuf_io_deq_valid),
    .io_deq_bits_listenAddr(cpu2_lbuf_io_deq_bits_listenAddr)
  );
  DFCExptArbiter expt_arbiter ( // @[DFCTable.scala 115:28]
    .io_table_e_data_ready(expt_arbiter_io_table_e_data_ready),
    .io_table_e_data_valid(expt_arbiter_io_table_e_data_valid),
    .io_table_e_data_bits_pid(expt_arbiter_io_table_e_data_bits_pid),
    .io_cpu1_e_data_ready(expt_arbiter_io_cpu1_e_data_ready),
    .io_cpu1_e_data_valid(expt_arbiter_io_cpu1_e_data_valid),
    .io_cpu1_e_data_bits_pid(expt_arbiter_io_cpu1_e_data_bits_pid)
  );
  assign io_cpu1_e_data_valid = expt_arbiter_io_cpu1_e_data_valid; // @[DFCTable.scala 137:13]
  assign io_cpu1_e_data_bits_pid = expt_arbiter_io_cpu1_e_data_bits_pid; // @[DFCTable.scala 137:13]
  assign io_cpu_f_data_valid = dfc_tableA_io_dfc_full_data_valid; // @[DFCTable.scala 141:12]
  assign io_cpu_f_data_bits_full_sig = dfc_tableA_io_dfc_full_data_bits_full_sig; // @[DFCTable.scala 141:12]
  assign dfc_tableA_clock = clock;
  assign dfc_tableA_reset = reset;
  assign dfc_tableA_io_cpu_w_data_valid = dfc_arbiter_io_table_w_data_valid; // @[DFCTable.scala 121:23]
  assign dfc_tableA_io_cpu_w_data_bits_listenAddr = dfc_arbiter_io_table_w_data_bits_listenAddr; // @[DFCTable.scala 121:23]
  assign dfc_tableA_io_cpu_w_data_bits_wPid = dfc_arbiter_io_table_w_data_bits_wPid; // @[DFCTable.scala 121:23]
  assign dfc_tableA_io_cpu_l_data_valid = dfc_arbiter_io_table_l_data_valid; // @[DFCTable.scala 122:23]
  assign dfc_tableA_io_cpu_l_data_bits_listenAddr = dfc_arbiter_io_table_l_data_bits_listenAddr; // @[DFCTable.scala 122:23]
  assign dfc_tableA_io_tableD_wdata_ready = dfc_tableD_io_tableA_wdata_ready; // @[DFCTable.scala 118:24]
  assign dfc_tableA_io_tableD_ldata_ready = dfc_tableD_io_tableA_ldata_ready; // @[DFCTable.scala 118:24]
  assign dfc_tableA_io_tableD_wresp_valid = dfc_tableD_io_tableA_wresp_valid; // @[DFCTable.scala 118:24]
  assign dfc_tableA_io_tableD_wresp_bits = dfc_tableD_io_tableA_wresp_bits; // @[DFCTable.scala 118:24]
  assign dfc_tableA_io_tableD_lresp_valid = dfc_tableD_io_tableA_lresp_valid; // @[DFCTable.scala 118:24]
  assign dfc_tableA_io_tableD_lresp_bits_tableAId = dfc_tableD_io_tableA_lresp_bits_tableAId; // @[DFCTable.scala 118:24]
  assign dfc_tableA_io_tableD_lresp_bits_finish = dfc_tableD_io_tableA_lresp_bits_finish; // @[DFCTable.scala 118:24]
  assign dfc_tableA_io_cpu_expt_data_ready = expt_arbiter_io_table_e_data_ready; // @[DFCTable.scala 139:27]
  assign dfc_tableD_clock = clock;
  assign dfc_tableD_reset = reset;
  assign dfc_tableD_io_tableA_wdata_valid = dfc_tableA_io_tableD_wdata_valid; // @[DFCTable.scala 118:24]
  assign dfc_tableD_io_tableA_wdata_bits_listenAddr = dfc_tableA_io_tableD_wdata_bits_listenAddr; // @[DFCTable.scala 118:24]
  assign dfc_tableD_io_tableA_wdata_bits_tableAId = dfc_tableA_io_tableD_wdata_bits_tableAId; // @[DFCTable.scala 118:24]
  assign dfc_tableD_io_tableA_ldata_valid = dfc_tableA_io_tableD_ldata_valid; // @[DFCTable.scala 118:24]
  assign dfc_tableD_io_tableA_ldata_bits_listenAddr = dfc_tableA_io_tableD_ldata_bits_listenAddr; // @[DFCTable.scala 118:24]
  assign dfc_tableD_io_tableA_wresp_ready = dfc_tableA_io_tableD_wresp_ready; // @[DFCTable.scala 118:24]
  assign dfc_tableD_io_tableA_lresp_ready = dfc_tableA_io_tableD_lresp_ready; // @[DFCTable.scala 118:24]
  assign dfc_arbiter_io_cpu1_w_data_valid = cpu1_wbuf_io_deq_valid; // @[DFCTable.scala 125:30]
  assign dfc_arbiter_io_cpu1_w_data_bits_listenAddr = cpu1_wbuf_io_deq_bits_listenAddr; // @[DFCTable.scala 125:30]
  assign dfc_arbiter_io_cpu1_w_data_bits_wPid = cpu1_wbuf_io_deq_bits_wPid; // @[DFCTable.scala 125:30]
  assign dfc_arbiter_io_cpu2_w_data_valid = cpu2_wbuf_io_deq_valid; // @[DFCTable.scala 127:30]
  assign dfc_arbiter_io_cpu2_w_data_bits_listenAddr = cpu2_wbuf_io_deq_bits_listenAddr; // @[DFCTable.scala 127:30]
  assign dfc_arbiter_io_cpu2_w_data_bits_wPid = cpu2_wbuf_io_deq_bits_wPid; // @[DFCTable.scala 127:30]
  assign dfc_arbiter_io_cpu1_l_data_valid = cpu1_lbuf_io_deq_valid; // @[DFCTable.scala 126:30]
  assign dfc_arbiter_io_cpu1_l_data_bits_listenAddr = cpu1_lbuf_io_deq_bits_listenAddr; // @[DFCTable.scala 126:30]
  assign dfc_arbiter_io_cpu2_l_data_valid = cpu2_lbuf_io_deq_valid; // @[DFCTable.scala 128:30]
  assign dfc_arbiter_io_cpu2_l_data_bits_listenAddr = cpu2_lbuf_io_deq_bits_listenAddr; // @[DFCTable.scala 128:30]
  assign dfc_arbiter_io_table_w_data_ready = dfc_tableA_io_cpu_w_data_ready; // @[DFCTable.scala 121:23]
  assign dfc_arbiter_io_table_l_data_ready = dfc_tableA_io_cpu_l_data_ready; // @[DFCTable.scala 122:23]
  assign cpu1_wbuf_clock = clock;
  assign cpu1_wbuf_reset = reset;
  assign cpu1_wbuf_io_enq_valid = io_cpu1_w_data_valid; // @[DFCTable.scala 131:20]
  assign cpu1_wbuf_io_enq_bits_listenAddr = io_cpu1_w_data_bits_listenAddr; // @[DFCTable.scala 131:20]
  assign cpu1_wbuf_io_enq_bits_wPid = io_cpu1_w_data_bits_wPid; // @[DFCTable.scala 131:20]
  assign cpu1_wbuf_io_deq_ready = dfc_arbiter_io_cpu1_w_data_ready; // @[DFCTable.scala 125:30]
  assign cpu2_wbuf_clock = clock;
  assign cpu2_wbuf_reset = reset;
  assign cpu2_wbuf_io_enq_valid = 1'h0; // @[DFCTable.scala 133:20]
  assign cpu2_wbuf_io_enq_bits_listenAddr = 32'h0; // @[DFCTable.scala 133:20]
  assign cpu2_wbuf_io_enq_bits_wPid = 16'h0; // @[DFCTable.scala 133:20]
  assign cpu2_wbuf_io_deq_ready = dfc_arbiter_io_cpu2_w_data_ready; // @[DFCTable.scala 127:30]
  assign cpu1_lbuf_clock = clock;
  assign cpu1_lbuf_reset = reset;
  assign cpu1_lbuf_io_enq_valid = io_cpu1_l_data_valid; // @[DFCTable.scala 132:20]
  assign cpu1_lbuf_io_enq_bits_listenAddr = io_cpu1_l_data_bits_listenAddr; // @[DFCTable.scala 132:20]
  assign cpu1_lbuf_io_deq_ready = dfc_arbiter_io_cpu1_l_data_ready; // @[DFCTable.scala 126:30]
  assign cpu2_lbuf_clock = clock;
  assign cpu2_lbuf_reset = reset;
  assign cpu2_lbuf_io_enq_valid = 1'h0; // @[DFCTable.scala 134:20]
  assign cpu2_lbuf_io_enq_bits_listenAddr = 32'h0; // @[DFCTable.scala 134:20]
  assign cpu2_lbuf_io_deq_ready = dfc_arbiter_io_cpu2_l_data_ready; // @[DFCTable.scala 128:30]
  assign expt_arbiter_io_table_e_data_valid = dfc_tableA_io_cpu_expt_data_valid; // @[DFCTable.scala 139:27]
  assign expt_arbiter_io_table_e_data_bits_pid = dfc_tableA_io_cpu_expt_data_bits_pid; // @[DFCTable.scala 139:27]
  assign expt_arbiter_io_cpu1_e_data_ready = io_cpu1_e_data_ready; // @[DFCTable.scala 137:13]
endmodule
module CSR(
  input         clock,
  input         reset,
  input         io__stall,
  input  [2:0]  io__cmd,
  input  [31:0] io__in,
  output [31:0] io__out,
  input  [31:0] io__pc,
  input  [31:0] io__addr,
  input  [31:0] io__inst,
  input         io__illegal,
  input  [1:0]  io__st_type,
  input  [2:0]  io__ld_type,
  input         io__pc_check,
  output        io__expt,
  output [31:0] io__evec,
  output [31:0] io__epc,
  output        io__vmSwitch,
  output [31:0] io__vmSwitchPC,
  input  [2:0]  io__dfc_cmd,
  input  [15:0] io__dfc_pid,
  input         io__table_f_data_valid,
  input         io__table_f_data_bits_full_sig,
  output        io__dfc_full,
  input         uartRxValid_0,
  input  [1:0]  dmmu,
  output        io_vmSwitch,
  output [31:0] io_in,
  output        clearPageFault_0,
  input  [1:0]  immu,
  output [31:0] satp_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire [11:0] csr_addr = io__inst[31:20]; // @[CSR.scala 128:25]
  wire [4:0] rs1_addr = io__inst[19:15]; // @[CSR.scala 129:25]
  reg [31:0] time_; // @[CSR.scala 132:25]
  reg [31:0] counter; // @[CSR.scala 133:25]
  reg [31:0] timeh; // @[CSR.scala 134:25]
  reg [31:0] cycle; // @[CSR.scala 135:25]
  reg [31:0] cycleh; // @[CSR.scala 136:25]
  reg [31:0] instret; // @[CSR.scala 137:25]
  reg [31:0] instreth; // @[CSR.scala 138:25]
  reg [1:0] PRV; // @[CSR.scala 147:21]
  reg [1:0] PRV1; // @[CSR.scala 148:21]
  reg  IE; // @[CSR.scala 151:20]
  reg  IE1; // @[CSR.scala 152:20]
  wire [31:0] mstatus = {22'h0,3'h0,1'h0,PRV1,IE1,PRV,IE}; // @[Cat.scala 30:58]
  reg [31:0] mtvec; // @[CSR.scala 164:24]
  reg  MTIP; // @[CSR.scala 168:21]
  reg  MTIE; // @[CSR.scala 171:21]
  reg  MSIP; // @[CSR.scala 174:21]
  reg  MSIE; // @[CSR.scala 177:21]
  wire [31:0] mip = {24'h0,MTIP,1'h0,2'h0,MSIP,1'h0,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] mie = {24'h0,MTIE,1'h0,2'h0,MSIE,1'h0,2'h0}; // @[Cat.scala 30:58]
  reg  uartInterruptPending; // @[CSR.scala 183:37]
  reg [31:0] mtimecmp; // @[CSR.scala 185:21]
  reg [31:0] mscratch; // @[CSR.scala 187:21]
  reg [31:0] mepc; // @[CSR.scala 189:17]
  reg [31:0] mcause; // @[CSR.scala 190:19]
  reg [31:0] mbadaddr; // @[CSR.scala 191:21]
  reg [31:0] mtohost; // @[CSR.scala 193:24]
  reg [31:0] mfromhost; // @[CSR.scala 194:22]
  reg [31:0] satp; // @[CSR.scala 202:21]
  wire [1:0] pageFault = immu != 2'h0 ? immu : dmmu; // @[CSR.scala 207:22]
  wire  _GEN_1 = uartRxValid_0 | uartInterruptPending; // @[CSR.scala 221:20 CSR.scala 221:42 CSR.scala 183:37]
  reg [31:0] dfc_pid; // @[CSR.scala 224:24]
  reg  dfc_full_reg; // @[CSR.scala 225:29]
  wire  _T_2 = 12'hc00 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_4 = 12'hc01 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_6 = 12'hc02 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_8 = 12'hc80 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_10 = 12'hc81 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_12 = 12'hc82 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_14 = 12'h900 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_16 = 12'h901 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_18 = 12'h902 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_20 = 12'h980 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_22 = 12'h981 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_24 = 12'h982 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_26 = 12'hf00 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_28 = 12'hf01 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_30 = 12'hf10 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_32 = 12'h301 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_34 = 12'h302 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_36 = 12'h304 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_38 = 12'h321 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_40 = 12'h701 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_42 = 12'h741 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_44 = 12'h340 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_46 = 12'h341 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_48 = 12'h342 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_50 = 12'h343 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_52 = 12'h344 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_54 = 12'h780 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_56 = 12'h781 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_58 = 12'h300 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_60 = 12'h180 == csr_addr; // @[Lookup.scala 31:38]
  wire  _T_62 = 12'h800 == csr_addr; // @[Lookup.scala 31:38]
  wire [31:0] _T_63 = _T_62 ? dfc_pid : 32'h0; // @[Lookup.scala 33:37]
  wire [31:0] _T_64 = _T_60 ? satp : _T_63; // @[Lookup.scala 33:37]
  wire [31:0] _T_65 = _T_58 ? mstatus : _T_64; // @[Lookup.scala 33:37]
  wire [31:0] _T_66 = _T_56 ? mfromhost : _T_65; // @[Lookup.scala 33:37]
  wire [31:0] _T_67 = _T_54 ? mtohost : _T_66; // @[Lookup.scala 33:37]
  wire [31:0] _T_68 = _T_52 ? mip : _T_67; // @[Lookup.scala 33:37]
  wire [31:0] _T_69 = _T_50 ? mbadaddr : _T_68; // @[Lookup.scala 33:37]
  wire [31:0] _T_70 = _T_48 ? mcause : _T_69; // @[Lookup.scala 33:37]
  wire [31:0] _T_71 = _T_46 ? mepc : _T_70; // @[Lookup.scala 33:37]
  wire [31:0] _T_72 = _T_44 ? mscratch : _T_71; // @[Lookup.scala 33:37]
  wire [31:0] _T_73 = _T_42 ? timeh : _T_72; // @[Lookup.scala 33:37]
  wire [31:0] _T_74 = _T_40 ? time_ : _T_73; // @[Lookup.scala 33:37]
  wire [31:0] _T_75 = _T_38 ? mtimecmp : _T_74; // @[Lookup.scala 33:37]
  wire [31:0] _T_76 = _T_36 ? mie : _T_75; // @[Lookup.scala 33:37]
  wire [31:0] _T_77 = _T_34 ? 32'h0 : _T_76; // @[Lookup.scala 33:37]
  wire [31:0] _T_78 = _T_32 ? mtvec : _T_77; // @[Lookup.scala 33:37]
  wire [31:0] _T_79 = _T_30 ? 32'h0 : _T_78; // @[Lookup.scala 33:37]
  wire [31:0] _T_80 = _T_28 ? 32'h0 : _T_79; // @[Lookup.scala 33:37]
  wire [31:0] _T_81 = _T_26 ? 32'h100100 : _T_80; // @[Lookup.scala 33:37]
  wire [31:0] _T_82 = _T_24 ? instreth : _T_81; // @[Lookup.scala 33:37]
  wire [31:0] _T_83 = _T_22 ? timeh : _T_82; // @[Lookup.scala 33:37]
  wire [31:0] _T_84 = _T_20 ? cycleh : _T_83; // @[Lookup.scala 33:37]
  wire [31:0] _T_85 = _T_18 ? instret : _T_84; // @[Lookup.scala 33:37]
  wire [31:0] _T_86 = _T_16 ? time_ : _T_85; // @[Lookup.scala 33:37]
  wire [31:0] _T_87 = _T_14 ? cycle : _T_86; // @[Lookup.scala 33:37]
  wire [31:0] _T_88 = _T_12 ? instreth : _T_87; // @[Lookup.scala 33:37]
  wire [31:0] _T_89 = _T_10 ? timeh : _T_88; // @[Lookup.scala 33:37]
  wire [31:0] _T_90 = _T_8 ? cycleh : _T_89; // @[Lookup.scala 33:37]
  wire [31:0] _T_91 = _T_6 ? instret : _T_90; // @[Lookup.scala 33:37]
  wire [31:0] _T_92 = _T_4 ? time_ : _T_91; // @[Lookup.scala 33:37]
  wire  privValid = csr_addr[9:8] <= PRV; // @[CSR.scala 265:34]
  wire  privInst = io__cmd == 3'h4; // @[CSR.scala 266:26]
  wire  _T_97 = privInst & ~csr_addr[0]; // @[CSR.scala 267:28]
  wire  _T_99 = ~csr_addr[8]; // @[CSR.scala 267:47]
  wire  isEcall = privInst & ~csr_addr[0] & ~csr_addr[8]; // @[CSR.scala 267:44]
  wire  isEbreak = privInst & csr_addr[0] & _T_99; // @[CSR.scala 268:44]
  wire  isEret = _T_97 & csr_addr[8]; // @[CSR.scala 269:44]
  wire  csrValid = _T_2 | _T_4 | _T_6 | _T_8 | _T_10 | _T_12 | _T_14 | _T_16 | _T_18 | _T_20 | _T_22 | _T_24 | _T_26 |
    _T_28 | _T_30 | _T_32 | _T_34 | _T_36 | _T_38 | _T_40 | _T_42 | _T_44 | _T_46 | _T_48 | _T_50 | _T_52 | _T_54 |
    _T_56 | _T_58 | _T_60 | _T_62; // @[CSR.scala 270:61]
  wire  csrRO = &csr_addr[11:10] | csr_addr == 12'h302; // @[CSR.scala 271:41]
  wire  wen = io__cmd == 3'h1 | io__cmd[1] & |rs1_addr; // @[CSR.scala 272:36]
  wire [31:0] _T_206 = io__out | io__in; // @[CSR.scala 275:22]
  wire [31:0] _T_207 = ~io__in; // @[CSR.scala 276:24]
  wire [31:0] _T_208 = io__out & _T_207; // @[CSR.scala 276:22]
  wire [31:0] _T_210 = 3'h1 == io__cmd ? io__in : 32'h0; // @[Mux.scala 80:57]
  wire [31:0] _T_212 = 3'h2 == io__cmd ? _T_206 : _T_210; // @[Mux.scala 80:57]
  wire [31:0] wdata = 3'h3 == io__cmd ? _T_208 : _T_212; // @[Mux.scala 80:57]
  wire  iaddrInvalid = io__pc_check & io__addr[1]; // @[CSR.scala 278:34]
  wire  _T_216 = |io__addr[1:0]; // @[CSR.scala 280:36]
  wire  _T_222 = 3'h2 == io__ld_type ? io__addr[0] : 3'h1 == io__ld_type & _T_216; // @[Mux.scala 80:57]
  wire  laddrInvalid = 3'h4 == io__ld_type ? io__addr[0] : _T_222; // @[Mux.scala 80:57]
  wire  saddrInvalid = 2'h2 == io__st_type ? io__addr[0] : 2'h1 == io__st_type & _T_216; // @[Mux.scala 80:57]
  wire  isInstructionFault = pageFault == 2'h1; // @[CSR.scala 284:38]
  wire  isLoadFault = pageFault == 2'h2; // @[CSR.scala 285:38]
  wire  isStoreFault = pageFault == 2'h3; // @[CSR.scala 286:38]
  wire  _T_230 = csr_addr == 12'h180; // @[CSR.scala 288:27]
  reg [31:0] vmSwitchPC; // @[CSR.scala 289:27]
  wire  _T_233 = io__inst != 32'h13; // @[CSR.scala 293:64]
  wire  _T_235 = pageFault == 2'h0; // @[CSR.scala 293:89]
  wire  isUartInterrupt = IE & uartInterruptPending & io__inst != 32'h13 & pageFault == 2'h0; // @[CSR.scala 293:86]
  wire  isTimerInterrupt = MTIP & MTIE & IE & _T_233 & _T_235 & ~isUartInterrupt; // @[CSR.scala 294:93]
  wire  isDFCAct = |io__dfc_pid; // @[CSR.scala 297:33]
  wire  writeDFCInvalid = dfc_full_reg & io__dfc_cmd == 3'h1; // @[CSR.scala 298:38]
  wire  _T_250 = ~privValid; // @[CSR.scala 306:51]
  wire  _T_252 = |io__cmd[1:0] & (~csrValid | ~privValid); // @[CSR.scala 306:34]
  wire  _T_253 = io__illegal | iaddrInvalid | laddrInvalid | saddrInvalid | _T_252; // @[CSR.scala 305:75]
  wire  _T_257 = privInst & _T_250; // @[CSR.scala 307:27]
  wire  _T_258 = _T_253 | wen & csrRO | _T_257; // @[CSR.scala 306:79]
  wire  _T_262 = _T_258 | isEcall | isEbreak | isInstructionFault | isLoadFault; // @[CSR.scala 307:86]
  wire  t_expt = _T_262 | isStoreFault | isTimerInterrupt | isUartInterrupt; // @[CSR.scala 308:65]
  wire [31:0] _T_268 = counter + 32'h1; // @[CSR.scala 315:22]
  wire [31:0] _T_272 = time_ + 32'h1; // @[CSR.scala 316:44]
  wire [31:0] _GEN_4 = &counter[10:0] ? _T_272 : time_; // @[CSR.scala 316:29 CSR.scala 316:36 CSR.scala 132:25]
  wire [31:0] _T_275 = timeh + 32'h1; // @[CSR.scala 317:36]
  wire [31:0] _GEN_5 = &time_ ? _T_275 : timeh; // @[CSR.scala 317:19 CSR.scala 317:27 CSR.scala 134:25]
  wire  _GEN_6 = time_ == mtimecmp | MTIP; // @[CSR.scala 318:26 CSR.scala 318:32 CSR.scala 168:21]
  wire [31:0] _T_278 = cycle + 32'h1; // @[CSR.scala 320:18]
  wire [31:0] _T_281 = cycleh + 32'h1; // @[CSR.scala 321:39]
  wire [31:0] _GEN_7 = &cycle ? _T_281 : cycleh; // @[CSR.scala 321:20 CSR.scala 321:29 CSR.scala 136:25]
  wire  _T_287 = ~io__stall; // @[CSR.scala 322:88]
  wire  isInstRet = _T_233 & (~io__expt | isEcall | isEbreak) & ~io__stall; // @[CSR.scala 322:85]
  wire [31:0] _T_289 = instret + 32'h1; // @[CSR.scala 323:40]
  wire [31:0] _GEN_8 = isInstRet ? _T_289 : instret; // @[CSR.scala 323:19 CSR.scala 323:29 CSR.scala 137:25]
  wire [31:0] _T_293 = instreth + 32'h1; // @[CSR.scala 324:58]
  wire [31:0] _GEN_9 = isInstRet & &instret ? _T_293 : instreth; // @[CSR.scala 324:35 CSR.scala 324:46 CSR.scala 138:25]
  wire [31:0] _T_296 = {io__pc[31:2], 2'h0}; // @[CSR.scala 328:28]
  wire [3:0] _GEN_345 = {{2'd0}, PRV}; // @[CSR.scala 335:47]
  wire [3:0] _T_298 = 4'h8 + _GEN_345; // @[CSR.scala 335:47]
  wire [4:0] _T_299 = writeDFCInvalid ? 5'h14 : 5'h2; // @[CSR.scala 346:20]
  wire [4:0] _T_300 = isUartInterrupt ? 5'h10 : _T_299; // @[CSR.scala 344:20]
  wire [31:0] _T_301 = isTimerInterrupt ? 32'h80000001 : {{27'd0}, _T_300}; // @[CSR.scala 342:20]
  wire [31:0] _T_302 = isStoreFault ? 32'hf : _T_301; // @[CSR.scala 340:20]
  wire [31:0] _T_303 = isLoadFault ? 32'hd : _T_302; // @[CSR.scala 339:20]
  wire [31:0] _T_304 = isInstructionFault ? 32'hc : _T_303; // @[CSR.scala 338:20]
  wire [31:0] _T_305 = isEbreak ? 32'h3 : _T_304; // @[CSR.scala 336:20]
  wire [31:0] _T_306 = isEcall ? {{28'd0}, _T_298} : _T_305; // @[CSR.scala 335:20]
  wire [31:0] _T_307 = saddrInvalid ? 32'h6 : _T_306; // @[CSR.scala 334:20]
  wire [31:0] _T_308 = laddrInvalid ? 32'h4 : _T_307; // @[CSR.scala 333:20]
  wire  _T_317 = isInstructionFault | isLoadFault | isStoreFault; // @[CSR.scala 354:46]
  wire [31:0] _T_326 = {{2'd0}, wdata[31:2]}; // @[CSR.scala 379:56]
  wire [33:0] _GEN_347 = {_T_326, 2'h0}; // @[CSR.scala 379:63]
  wire [34:0] _T_327 = {{1'd0}, _GEN_347}; // @[CSR.scala 379:63]
  wire [31:0] _GEN_13 = csr_addr == 12'h301 ? wdata : mtvec; // @[CSR.scala 392:41 CSR.scala 392:49 CSR.scala 164:24]
  wire [31:0] _GEN_14 = _T_230 ? wdata : satp; // @[CSR.scala 391:40 CSR.scala 391:47 CSR.scala 202:21]
  wire [31:0] _GEN_15 = _T_230 ? io__pc : vmSwitchPC; // @[CSR.scala 391:40 CSR.scala 391:69 CSR.scala 289:27]
  wire [31:0] _GEN_16 = _T_230 ? mtvec : _GEN_13; // @[CSR.scala 391:40 CSR.scala 164:24]
  wire [31:0] _GEN_17 = csr_addr == 12'h982 ? wdata : _GEN_9; // @[CSR.scala 390:45 CSR.scala 390:56]
  wire [31:0] _GEN_18 = csr_addr == 12'h982 ? satp : _GEN_14; // @[CSR.scala 390:45 CSR.scala 202:21]
  wire [31:0] _GEN_19 = csr_addr == 12'h982 ? vmSwitchPC : _GEN_15; // @[CSR.scala 390:45 CSR.scala 289:27]
  wire [31:0] _GEN_20 = csr_addr == 12'h982 ? mtvec : _GEN_16; // @[CSR.scala 390:45 CSR.scala 164:24]
  wire [31:0] _GEN_21 = csr_addr == 12'h981 ? wdata : _GEN_5; // @[CSR.scala 389:42 CSR.scala 389:50]
  wire [31:0] _GEN_22 = csr_addr == 12'h981 ? _GEN_9 : _GEN_17; // @[CSR.scala 389:42]
  wire [31:0] _GEN_23 = csr_addr == 12'h981 ? satp : _GEN_18; // @[CSR.scala 389:42 CSR.scala 202:21]
  wire [31:0] _GEN_24 = csr_addr == 12'h981 ? vmSwitchPC : _GEN_19; // @[CSR.scala 389:42 CSR.scala 289:27]
  wire [31:0] _GEN_25 = csr_addr == 12'h981 ? mtvec : _GEN_20; // @[CSR.scala 389:42 CSR.scala 164:24]
  wire [31:0] _GEN_26 = csr_addr == 12'h980 ? wdata : _GEN_7; // @[CSR.scala 388:43 CSR.scala 388:52]
  wire [31:0] _GEN_27 = csr_addr == 12'h980 ? _GEN_5 : _GEN_21; // @[CSR.scala 388:43]
  wire [31:0] _GEN_28 = csr_addr == 12'h980 ? _GEN_9 : _GEN_22; // @[CSR.scala 388:43]
  wire [31:0] _GEN_29 = csr_addr == 12'h980 ? satp : _GEN_23; // @[CSR.scala 388:43 CSR.scala 202:21]
  wire [31:0] _GEN_30 = csr_addr == 12'h980 ? vmSwitchPC : _GEN_24; // @[CSR.scala 388:43 CSR.scala 289:27]
  wire [31:0] _GEN_31 = csr_addr == 12'h980 ? mtvec : _GEN_25; // @[CSR.scala 388:43 CSR.scala 164:24]
  wire [31:0] _GEN_32 = csr_addr == 12'h902 ? wdata : _GEN_8; // @[CSR.scala 387:44 CSR.scala 387:54]
  wire [31:0] _GEN_33 = csr_addr == 12'h902 ? _GEN_7 : _GEN_26; // @[CSR.scala 387:44]
  wire [31:0] _GEN_34 = csr_addr == 12'h902 ? _GEN_5 : _GEN_27; // @[CSR.scala 387:44]
  wire [31:0] _GEN_35 = csr_addr == 12'h902 ? _GEN_9 : _GEN_28; // @[CSR.scala 387:44]
  wire [31:0] _GEN_36 = csr_addr == 12'h902 ? satp : _GEN_29; // @[CSR.scala 387:44 CSR.scala 202:21]
  wire [31:0] _GEN_37 = csr_addr == 12'h902 ? vmSwitchPC : _GEN_30; // @[CSR.scala 387:44 CSR.scala 289:27]
  wire [31:0] _GEN_38 = csr_addr == 12'h902 ? mtvec : _GEN_31; // @[CSR.scala 387:44 CSR.scala 164:24]
  wire [31:0] _GEN_39 = csr_addr == 12'h901 ? wdata : _GEN_4; // @[CSR.scala 386:41 CSR.scala 386:48]
  wire [31:0] _GEN_40 = csr_addr == 12'h901 ? _GEN_8 : _GEN_32; // @[CSR.scala 386:41]
  wire [31:0] _GEN_41 = csr_addr == 12'h901 ? _GEN_7 : _GEN_33; // @[CSR.scala 386:41]
  wire [31:0] _GEN_42 = csr_addr == 12'h901 ? _GEN_5 : _GEN_34; // @[CSR.scala 386:41]
  wire [31:0] _GEN_43 = csr_addr == 12'h901 ? _GEN_9 : _GEN_35; // @[CSR.scala 386:41]
  wire [31:0] _GEN_44 = csr_addr == 12'h901 ? satp : _GEN_36; // @[CSR.scala 386:41 CSR.scala 202:21]
  wire [31:0] _GEN_45 = csr_addr == 12'h901 ? vmSwitchPC : _GEN_37; // @[CSR.scala 386:41 CSR.scala 289:27]
  wire [31:0] _GEN_46 = csr_addr == 12'h901 ? mtvec : _GEN_38; // @[CSR.scala 386:41 CSR.scala 164:24]
  wire [31:0] _GEN_47 = csr_addr == 12'h900 ? wdata : _T_278; // @[CSR.scala 385:42 CSR.scala 385:50 CSR.scala 320:9]
  wire [31:0] _GEN_48 = csr_addr == 12'h900 ? _GEN_4 : _GEN_39; // @[CSR.scala 385:42]
  wire [31:0] _GEN_49 = csr_addr == 12'h900 ? _GEN_8 : _GEN_40; // @[CSR.scala 385:42]
  wire [31:0] _GEN_50 = csr_addr == 12'h900 ? _GEN_7 : _GEN_41; // @[CSR.scala 385:42]
  wire [31:0] _GEN_51 = csr_addr == 12'h900 ? _GEN_5 : _GEN_42; // @[CSR.scala 385:42]
  wire [31:0] _GEN_52 = csr_addr == 12'h900 ? _GEN_9 : _GEN_43; // @[CSR.scala 385:42]
  wire [31:0] _GEN_53 = csr_addr == 12'h900 ? satp : _GEN_44; // @[CSR.scala 385:42 CSR.scala 202:21]
  wire [31:0] _GEN_54 = csr_addr == 12'h900 ? vmSwitchPC : _GEN_45; // @[CSR.scala 385:42 CSR.scala 289:27]
  wire [31:0] _GEN_55 = csr_addr == 12'h900 ? mtvec : _GEN_46; // @[CSR.scala 385:42 CSR.scala 164:24]
  wire [31:0] _GEN_56 = csr_addr == 12'h781 ? wdata : mfromhost; // @[CSR.scala 384:45 CSR.scala 384:57]
  wire [31:0] _GEN_57 = csr_addr == 12'h781 ? _T_278 : _GEN_47; // @[CSR.scala 384:45 CSR.scala 320:9]
  wire [31:0] _GEN_58 = csr_addr == 12'h781 ? _GEN_4 : _GEN_48; // @[CSR.scala 384:45]
  wire [31:0] _GEN_59 = csr_addr == 12'h781 ? _GEN_8 : _GEN_49; // @[CSR.scala 384:45]
  wire [31:0] _GEN_60 = csr_addr == 12'h781 ? _GEN_7 : _GEN_50; // @[CSR.scala 384:45]
  wire [31:0] _GEN_61 = csr_addr == 12'h781 ? _GEN_5 : _GEN_51; // @[CSR.scala 384:45]
  wire [31:0] _GEN_62 = csr_addr == 12'h781 ? _GEN_9 : _GEN_52; // @[CSR.scala 384:45]
  wire [31:0] _GEN_63 = csr_addr == 12'h781 ? satp : _GEN_53; // @[CSR.scala 384:45 CSR.scala 202:21]
  wire [31:0] _GEN_64 = csr_addr == 12'h781 ? vmSwitchPC : _GEN_54; // @[CSR.scala 384:45 CSR.scala 289:27]
  wire [31:0] _GEN_65 = csr_addr == 12'h781 ? mtvec : _GEN_55; // @[CSR.scala 384:45 CSR.scala 164:24]
  wire [31:0] _GEN_66 = csr_addr == 12'h780 ? wdata : mtohost; // @[CSR.scala 383:43 CSR.scala 383:53 CSR.scala 193:24]
  wire [31:0] _GEN_67 = csr_addr == 12'h780 ? mfromhost : _GEN_56; // @[CSR.scala 383:43]
  wire [31:0] _GEN_68 = csr_addr == 12'h780 ? _T_278 : _GEN_57; // @[CSR.scala 383:43 CSR.scala 320:9]
  wire [31:0] _GEN_69 = csr_addr == 12'h780 ? _GEN_4 : _GEN_58; // @[CSR.scala 383:43]
  wire [31:0] _GEN_70 = csr_addr == 12'h780 ? _GEN_8 : _GEN_59; // @[CSR.scala 383:43]
  wire [31:0] _GEN_71 = csr_addr == 12'h780 ? _GEN_7 : _GEN_60; // @[CSR.scala 383:43]
  wire [31:0] _GEN_72 = csr_addr == 12'h780 ? _GEN_5 : _GEN_61; // @[CSR.scala 383:43]
  wire [31:0] _GEN_73 = csr_addr == 12'h780 ? _GEN_9 : _GEN_62; // @[CSR.scala 383:43]
  wire [31:0] _GEN_74 = csr_addr == 12'h780 ? satp : _GEN_63; // @[CSR.scala 383:43 CSR.scala 202:21]
  wire [31:0] _GEN_75 = csr_addr == 12'h780 ? vmSwitchPC : _GEN_64; // @[CSR.scala 383:43 CSR.scala 289:27]
  wire [31:0] _GEN_76 = csr_addr == 12'h780 ? mtvec : _GEN_65; // @[CSR.scala 383:43 CSR.scala 164:24]
  wire [31:0] _GEN_77 = csr_addr == 12'h343 ? wdata : mbadaddr; // @[CSR.scala 382:44 CSR.scala 382:55 CSR.scala 191:21]
  wire [31:0] _GEN_78 = csr_addr == 12'h343 ? mtohost : _GEN_66; // @[CSR.scala 382:44 CSR.scala 193:24]
  wire [31:0] _GEN_79 = csr_addr == 12'h343 ? mfromhost : _GEN_67; // @[CSR.scala 382:44]
  wire [31:0] _GEN_80 = csr_addr == 12'h343 ? _T_278 : _GEN_68; // @[CSR.scala 382:44 CSR.scala 320:9]
  wire [31:0] _GEN_81 = csr_addr == 12'h343 ? _GEN_4 : _GEN_69; // @[CSR.scala 382:44]
  wire [31:0] _GEN_82 = csr_addr == 12'h343 ? _GEN_8 : _GEN_70; // @[CSR.scala 382:44]
  wire [31:0] _GEN_83 = csr_addr == 12'h343 ? _GEN_7 : _GEN_71; // @[CSR.scala 382:44]
  wire [31:0] _GEN_84 = csr_addr == 12'h343 ? _GEN_5 : _GEN_72; // @[CSR.scala 382:44]
  wire [31:0] _GEN_85 = csr_addr == 12'h343 ? _GEN_9 : _GEN_73; // @[CSR.scala 382:44]
  wire [31:0] _GEN_86 = csr_addr == 12'h343 ? satp : _GEN_74; // @[CSR.scala 382:44 CSR.scala 202:21]
  wire [31:0] _GEN_87 = csr_addr == 12'h343 ? vmSwitchPC : _GEN_75; // @[CSR.scala 382:44 CSR.scala 289:27]
  wire [31:0] _GEN_88 = csr_addr == 12'h343 ? mtvec : _GEN_76; // @[CSR.scala 382:44 CSR.scala 164:24]
  wire [31:0] _GEN_89 = csr_addr == 12'h342 ? wdata : mcause; // @[CSR.scala 381:42 CSR.scala 381:51 CSR.scala 190:19]
  wire [31:0] _GEN_90 = csr_addr == 12'h342 ? mbadaddr : _GEN_77; // @[CSR.scala 381:42 CSR.scala 191:21]
  wire [31:0] _GEN_91 = csr_addr == 12'h342 ? mtohost : _GEN_78; // @[CSR.scala 381:42 CSR.scala 193:24]
  wire [31:0] _GEN_92 = csr_addr == 12'h342 ? mfromhost : _GEN_79; // @[CSR.scala 381:42]
  wire [31:0] _GEN_93 = csr_addr == 12'h342 ? _T_278 : _GEN_80; // @[CSR.scala 381:42 CSR.scala 320:9]
  wire [31:0] _GEN_94 = csr_addr == 12'h342 ? _GEN_4 : _GEN_81; // @[CSR.scala 381:42]
  wire [31:0] _GEN_95 = csr_addr == 12'h342 ? _GEN_8 : _GEN_82; // @[CSR.scala 381:42]
  wire [31:0] _GEN_96 = csr_addr == 12'h342 ? _GEN_7 : _GEN_83; // @[CSR.scala 381:42]
  wire [31:0] _GEN_97 = csr_addr == 12'h342 ? _GEN_5 : _GEN_84; // @[CSR.scala 381:42]
  wire [31:0] _GEN_98 = csr_addr == 12'h342 ? _GEN_9 : _GEN_85; // @[CSR.scala 381:42]
  wire [31:0] _GEN_99 = csr_addr == 12'h342 ? satp : _GEN_86; // @[CSR.scala 381:42 CSR.scala 202:21]
  wire [31:0] _GEN_100 = csr_addr == 12'h342 ? vmSwitchPC : _GEN_87; // @[CSR.scala 381:42 CSR.scala 289:27]
  wire [31:0] _GEN_101 = csr_addr == 12'h342 ? mtvec : _GEN_88; // @[CSR.scala 381:42 CSR.scala 164:24]
  wire [34:0] _GEN_102 = csr_addr == 12'h341 ? _T_327 : {{3'd0}, mepc}; // @[CSR.scala 379:40 CSR.scala 379:47 CSR.scala 189:17]
  wire [31:0] _GEN_103 = csr_addr == 12'h341 ? mcause : _GEN_89; // @[CSR.scala 379:40 CSR.scala 190:19]
  wire [31:0] _GEN_104 = csr_addr == 12'h341 ? mbadaddr : _GEN_90; // @[CSR.scala 379:40 CSR.scala 191:21]
  wire [31:0] _GEN_105 = csr_addr == 12'h341 ? mtohost : _GEN_91; // @[CSR.scala 379:40 CSR.scala 193:24]
  wire [31:0] _GEN_106 = csr_addr == 12'h341 ? mfromhost : _GEN_92; // @[CSR.scala 379:40]
  wire [31:0] _GEN_107 = csr_addr == 12'h341 ? _T_278 : _GEN_93; // @[CSR.scala 379:40 CSR.scala 320:9]
  wire [31:0] _GEN_108 = csr_addr == 12'h341 ? _GEN_4 : _GEN_94; // @[CSR.scala 379:40]
  wire [31:0] _GEN_109 = csr_addr == 12'h341 ? _GEN_8 : _GEN_95; // @[CSR.scala 379:40]
  wire [31:0] _GEN_110 = csr_addr == 12'h341 ? _GEN_7 : _GEN_96; // @[CSR.scala 379:40]
  wire [31:0] _GEN_111 = csr_addr == 12'h341 ? _GEN_5 : _GEN_97; // @[CSR.scala 379:40]
  wire [31:0] _GEN_112 = csr_addr == 12'h341 ? _GEN_9 : _GEN_98; // @[CSR.scala 379:40]
  wire [31:0] _GEN_113 = csr_addr == 12'h341 ? satp : _GEN_99; // @[CSR.scala 379:40 CSR.scala 202:21]
  wire [31:0] _GEN_114 = csr_addr == 12'h341 ? vmSwitchPC : _GEN_100; // @[CSR.scala 379:40 CSR.scala 289:27]
  wire [31:0] _GEN_115 = csr_addr == 12'h341 ? mtvec : _GEN_101; // @[CSR.scala 379:40 CSR.scala 164:24]
  wire [31:0] _GEN_116 = csr_addr == 12'h340 ? wdata : mscratch; // @[CSR.scala 378:44 CSR.scala 378:55 CSR.scala 187:21]
  wire [34:0] _GEN_117 = csr_addr == 12'h340 ? {{3'd0}, mepc} : _GEN_102; // @[CSR.scala 378:44 CSR.scala 189:17]
  wire [31:0] _GEN_118 = csr_addr == 12'h340 ? mcause : _GEN_103; // @[CSR.scala 378:44 CSR.scala 190:19]
  wire [31:0] _GEN_119 = csr_addr == 12'h340 ? mbadaddr : _GEN_104; // @[CSR.scala 378:44 CSR.scala 191:21]
  wire [31:0] _GEN_120 = csr_addr == 12'h340 ? mtohost : _GEN_105; // @[CSR.scala 378:44 CSR.scala 193:24]
  wire [31:0] _GEN_121 = csr_addr == 12'h340 ? mfromhost : _GEN_106; // @[CSR.scala 378:44]
  wire [31:0] _GEN_122 = csr_addr == 12'h340 ? _T_278 : _GEN_107; // @[CSR.scala 378:44 CSR.scala 320:9]
  wire [31:0] _GEN_123 = csr_addr == 12'h340 ? _GEN_4 : _GEN_108; // @[CSR.scala 378:44]
  wire [31:0] _GEN_124 = csr_addr == 12'h340 ? _GEN_8 : _GEN_109; // @[CSR.scala 378:44]
  wire [31:0] _GEN_125 = csr_addr == 12'h340 ? _GEN_7 : _GEN_110; // @[CSR.scala 378:44]
  wire [31:0] _GEN_126 = csr_addr == 12'h340 ? _GEN_5 : _GEN_111; // @[CSR.scala 378:44]
  wire [31:0] _GEN_127 = csr_addr == 12'h340 ? _GEN_9 : _GEN_112; // @[CSR.scala 378:44]
  wire [31:0] _GEN_128 = csr_addr == 12'h340 ? satp : _GEN_113; // @[CSR.scala 378:44 CSR.scala 202:21]
  wire [31:0] _GEN_129 = csr_addr == 12'h340 ? vmSwitchPC : _GEN_114; // @[CSR.scala 378:44 CSR.scala 289:27]
  wire [31:0] _GEN_130 = csr_addr == 12'h340 ? mtvec : _GEN_115; // @[CSR.scala 378:44 CSR.scala 164:24]
  wire [31:0] _GEN_131 = csr_addr == 12'h321 ? wdata : mtimecmp; // @[CSR.scala 377:44 CSR.scala 377:55 CSR.scala 185:21]
  wire  _GEN_132 = csr_addr == 12'h321 ? 1'h0 : _GEN_6; // @[CSR.scala 377:44 CSR.scala 377:71]
  wire [31:0] _GEN_133 = csr_addr == 12'h321 ? mscratch : _GEN_116; // @[CSR.scala 377:44 CSR.scala 187:21]
  wire [34:0] _GEN_134 = csr_addr == 12'h321 ? {{3'd0}, mepc} : _GEN_117; // @[CSR.scala 377:44 CSR.scala 189:17]
  wire [31:0] _GEN_135 = csr_addr == 12'h321 ? mcause : _GEN_118; // @[CSR.scala 377:44 CSR.scala 190:19]
  wire [31:0] _GEN_136 = csr_addr == 12'h321 ? mbadaddr : _GEN_119; // @[CSR.scala 377:44 CSR.scala 191:21]
  wire [31:0] _GEN_137 = csr_addr == 12'h321 ? mtohost : _GEN_120; // @[CSR.scala 377:44 CSR.scala 193:24]
  wire [31:0] _GEN_138 = csr_addr == 12'h321 ? mfromhost : _GEN_121; // @[CSR.scala 377:44]
  wire [31:0] _GEN_139 = csr_addr == 12'h321 ? _T_278 : _GEN_122; // @[CSR.scala 377:44 CSR.scala 320:9]
  wire [31:0] _GEN_140 = csr_addr == 12'h321 ? _GEN_4 : _GEN_123; // @[CSR.scala 377:44]
  wire [31:0] _GEN_141 = csr_addr == 12'h321 ? _GEN_8 : _GEN_124; // @[CSR.scala 377:44]
  wire [31:0] _GEN_142 = csr_addr == 12'h321 ? _GEN_7 : _GEN_125; // @[CSR.scala 377:44]
  wire [31:0] _GEN_143 = csr_addr == 12'h321 ? _GEN_5 : _GEN_126; // @[CSR.scala 377:44]
  wire [31:0] _GEN_144 = csr_addr == 12'h321 ? _GEN_9 : _GEN_127; // @[CSR.scala 377:44]
  wire [31:0] _GEN_145 = csr_addr == 12'h321 ? satp : _GEN_128; // @[CSR.scala 377:44 CSR.scala 202:21]
  wire [31:0] _GEN_146 = csr_addr == 12'h321 ? vmSwitchPC : _GEN_129; // @[CSR.scala 377:44 CSR.scala 289:27]
  wire [31:0] _GEN_147 = csr_addr == 12'h321 ? mtvec : _GEN_130; // @[CSR.scala 377:44 CSR.scala 164:24]
  wire [31:0] _GEN_148 = csr_addr == 12'h741 ? wdata : _GEN_143; // @[CSR.scala 376:42 CSR.scala 376:50]
  wire [31:0] _GEN_149 = csr_addr == 12'h741 ? mtimecmp : _GEN_131; // @[CSR.scala 376:42 CSR.scala 185:21]
  wire  _GEN_150 = csr_addr == 12'h741 ? _GEN_6 : _GEN_132; // @[CSR.scala 376:42]
  wire [31:0] _GEN_151 = csr_addr == 12'h741 ? mscratch : _GEN_133; // @[CSR.scala 376:42 CSR.scala 187:21]
  wire [34:0] _GEN_152 = csr_addr == 12'h741 ? {{3'd0}, mepc} : _GEN_134; // @[CSR.scala 376:42 CSR.scala 189:17]
  wire [31:0] _GEN_153 = csr_addr == 12'h741 ? mcause : _GEN_135; // @[CSR.scala 376:42 CSR.scala 190:19]
  wire [31:0] _GEN_154 = csr_addr == 12'h741 ? mbadaddr : _GEN_136; // @[CSR.scala 376:42 CSR.scala 191:21]
  wire [31:0] _GEN_155 = csr_addr == 12'h741 ? mtohost : _GEN_137; // @[CSR.scala 376:42 CSR.scala 193:24]
  wire [31:0] _GEN_156 = csr_addr == 12'h741 ? mfromhost : _GEN_138; // @[CSR.scala 376:42]
  wire [31:0] _GEN_157 = csr_addr == 12'h741 ? _T_278 : _GEN_139; // @[CSR.scala 376:42 CSR.scala 320:9]
  wire [31:0] _GEN_158 = csr_addr == 12'h741 ? _GEN_4 : _GEN_140; // @[CSR.scala 376:42]
  wire [31:0] _GEN_159 = csr_addr == 12'h741 ? _GEN_8 : _GEN_141; // @[CSR.scala 376:42]
  wire [31:0] _GEN_160 = csr_addr == 12'h741 ? _GEN_7 : _GEN_142; // @[CSR.scala 376:42]
  wire [31:0] _GEN_161 = csr_addr == 12'h741 ? _GEN_9 : _GEN_144; // @[CSR.scala 376:42]
  wire [31:0] _GEN_162 = csr_addr == 12'h741 ? satp : _GEN_145; // @[CSR.scala 376:42 CSR.scala 202:21]
  wire [31:0] _GEN_163 = csr_addr == 12'h741 ? vmSwitchPC : _GEN_146; // @[CSR.scala 376:42 CSR.scala 289:27]
  wire [31:0] _GEN_164 = csr_addr == 12'h741 ? mtvec : _GEN_147; // @[CSR.scala 376:42 CSR.scala 164:24]
  wire [31:0] _GEN_165 = csr_addr == 12'h701 ? wdata : _GEN_158; // @[CSR.scala 375:41 CSR.scala 375:48]
  wire [31:0] _GEN_166 = csr_addr == 12'h701 ? _GEN_5 : _GEN_148; // @[CSR.scala 375:41]
  wire [31:0] _GEN_167 = csr_addr == 12'h701 ? mtimecmp : _GEN_149; // @[CSR.scala 375:41 CSR.scala 185:21]
  wire  _GEN_168 = csr_addr == 12'h701 ? _GEN_6 : _GEN_150; // @[CSR.scala 375:41]
  wire [31:0] _GEN_169 = csr_addr == 12'h701 ? mscratch : _GEN_151; // @[CSR.scala 375:41 CSR.scala 187:21]
  wire [34:0] _GEN_170 = csr_addr == 12'h701 ? {{3'd0}, mepc} : _GEN_152; // @[CSR.scala 375:41 CSR.scala 189:17]
  wire [31:0] _GEN_171 = csr_addr == 12'h701 ? mcause : _GEN_153; // @[CSR.scala 375:41 CSR.scala 190:19]
  wire [31:0] _GEN_172 = csr_addr == 12'h701 ? mbadaddr : _GEN_154; // @[CSR.scala 375:41 CSR.scala 191:21]
  wire [31:0] _GEN_173 = csr_addr == 12'h701 ? mtohost : _GEN_155; // @[CSR.scala 375:41 CSR.scala 193:24]
  wire [31:0] _GEN_174 = csr_addr == 12'h701 ? mfromhost : _GEN_156; // @[CSR.scala 375:41]
  wire [31:0] _GEN_175 = csr_addr == 12'h701 ? _T_278 : _GEN_157; // @[CSR.scala 375:41 CSR.scala 320:9]
  wire [31:0] _GEN_176 = csr_addr == 12'h701 ? _GEN_8 : _GEN_159; // @[CSR.scala 375:41]
  wire [31:0] _GEN_177 = csr_addr == 12'h701 ? _GEN_7 : _GEN_160; // @[CSR.scala 375:41]
  wire [31:0] _GEN_178 = csr_addr == 12'h701 ? _GEN_9 : _GEN_161; // @[CSR.scala 375:41]
  wire [31:0] _GEN_179 = csr_addr == 12'h701 ? satp : _GEN_162; // @[CSR.scala 375:41 CSR.scala 202:21]
  wire [31:0] _GEN_180 = csr_addr == 12'h701 ? vmSwitchPC : _GEN_163; // @[CSR.scala 375:41 CSR.scala 289:27]
  wire [31:0] _GEN_181 = csr_addr == 12'h701 ? mtvec : _GEN_164; // @[CSR.scala 375:41 CSR.scala 164:24]
  wire  _GEN_182 = csr_addr == 12'h304 ? wdata[7] : MTIE; // @[CSR.scala 371:39 CSR.scala 372:14 CSR.scala 171:21]
  wire  _GEN_183 = csr_addr == 12'h304 ? wdata[3] : MSIE; // @[CSR.scala 371:39 CSR.scala 373:14 CSR.scala 177:21]
  wire [31:0] _GEN_184 = csr_addr == 12'h304 ? _GEN_4 : _GEN_165; // @[CSR.scala 371:39]
  wire [31:0] _GEN_185 = csr_addr == 12'h304 ? _GEN_5 : _GEN_166; // @[CSR.scala 371:39]
  wire [31:0] _GEN_186 = csr_addr == 12'h304 ? mtimecmp : _GEN_167; // @[CSR.scala 371:39 CSR.scala 185:21]
  wire  _GEN_187 = csr_addr == 12'h304 ? _GEN_6 : _GEN_168; // @[CSR.scala 371:39]
  wire [31:0] _GEN_188 = csr_addr == 12'h304 ? mscratch : _GEN_169; // @[CSR.scala 371:39 CSR.scala 187:21]
  wire [34:0] _GEN_189 = csr_addr == 12'h304 ? {{3'd0}, mepc} : _GEN_170; // @[CSR.scala 371:39 CSR.scala 189:17]
  wire [31:0] _GEN_190 = csr_addr == 12'h304 ? mcause : _GEN_171; // @[CSR.scala 371:39 CSR.scala 190:19]
  wire [31:0] _GEN_191 = csr_addr == 12'h304 ? mbadaddr : _GEN_172; // @[CSR.scala 371:39 CSR.scala 191:21]
  wire [31:0] _GEN_192 = csr_addr == 12'h304 ? mtohost : _GEN_173; // @[CSR.scala 371:39 CSR.scala 193:24]
  wire [31:0] _GEN_193 = csr_addr == 12'h304 ? mfromhost : _GEN_174; // @[CSR.scala 371:39]
  wire [31:0] _GEN_194 = csr_addr == 12'h304 ? _T_278 : _GEN_175; // @[CSR.scala 371:39 CSR.scala 320:9]
  wire [31:0] _GEN_195 = csr_addr == 12'h304 ? _GEN_8 : _GEN_176; // @[CSR.scala 371:39]
  wire [31:0] _GEN_196 = csr_addr == 12'h304 ? _GEN_7 : _GEN_177; // @[CSR.scala 371:39]
  wire [31:0] _GEN_197 = csr_addr == 12'h304 ? _GEN_9 : _GEN_178; // @[CSR.scala 371:39]
  wire [31:0] _GEN_198 = csr_addr == 12'h304 ? satp : _GEN_179; // @[CSR.scala 371:39 CSR.scala 202:21]
  wire [31:0] _GEN_199 = csr_addr == 12'h304 ? vmSwitchPC : _GEN_180; // @[CSR.scala 371:39 CSR.scala 289:27]
  wire [31:0] _GEN_200 = csr_addr == 12'h304 ? mtvec : _GEN_181; // @[CSR.scala 371:39 CSR.scala 164:24]
  wire  _GEN_201 = csr_addr == 12'h344 ? wdata[7] : _GEN_187; // @[CSR.scala 367:39 CSR.scala 368:14]
  wire  _GEN_202 = csr_addr == 12'h344 ? wdata[3] : MSIP; // @[CSR.scala 367:39 CSR.scala 369:14 CSR.scala 174:21]
  wire  _GEN_203 = csr_addr == 12'h344 ? MTIE : _GEN_182; // @[CSR.scala 367:39 CSR.scala 171:21]
  wire  _GEN_204 = csr_addr == 12'h344 ? MSIE : _GEN_183; // @[CSR.scala 367:39 CSR.scala 177:21]
  wire [31:0] _GEN_205 = csr_addr == 12'h344 ? _GEN_4 : _GEN_184; // @[CSR.scala 367:39]
  wire [31:0] _GEN_206 = csr_addr == 12'h344 ? _GEN_5 : _GEN_185; // @[CSR.scala 367:39]
  wire [31:0] _GEN_207 = csr_addr == 12'h344 ? mtimecmp : _GEN_186; // @[CSR.scala 367:39 CSR.scala 185:21]
  wire [31:0] _GEN_208 = csr_addr == 12'h344 ? mscratch : _GEN_188; // @[CSR.scala 367:39 CSR.scala 187:21]
  wire [34:0] _GEN_209 = csr_addr == 12'h344 ? {{3'd0}, mepc} : _GEN_189; // @[CSR.scala 367:39 CSR.scala 189:17]
  wire [31:0] _GEN_210 = csr_addr == 12'h344 ? mcause : _GEN_190; // @[CSR.scala 367:39 CSR.scala 190:19]
  wire [31:0] _GEN_211 = csr_addr == 12'h344 ? mbadaddr : _GEN_191; // @[CSR.scala 367:39 CSR.scala 191:21]
  wire [31:0] _GEN_212 = csr_addr == 12'h344 ? mtohost : _GEN_192; // @[CSR.scala 367:39 CSR.scala 193:24]
  wire [31:0] _GEN_213 = csr_addr == 12'h344 ? mfromhost : _GEN_193; // @[CSR.scala 367:39]
  wire [31:0] _GEN_214 = csr_addr == 12'h344 ? _T_278 : _GEN_194; // @[CSR.scala 367:39 CSR.scala 320:9]
  wire [31:0] _GEN_215 = csr_addr == 12'h344 ? _GEN_8 : _GEN_195; // @[CSR.scala 367:39]
  wire [31:0] _GEN_216 = csr_addr == 12'h344 ? _GEN_7 : _GEN_196; // @[CSR.scala 367:39]
  wire [31:0] _GEN_217 = csr_addr == 12'h344 ? _GEN_9 : _GEN_197; // @[CSR.scala 367:39]
  wire [31:0] _GEN_218 = csr_addr == 12'h344 ? satp : _GEN_198; // @[CSR.scala 367:39 CSR.scala 202:21]
  wire [31:0] _GEN_219 = csr_addr == 12'h344 ? vmSwitchPC : _GEN_199; // @[CSR.scala 367:39 CSR.scala 289:27]
  wire [31:0] _GEN_220 = csr_addr == 12'h344 ? mtvec : _GEN_200; // @[CSR.scala 367:39 CSR.scala 164:24]
  wire [1:0] _GEN_221 = csr_addr == 12'h300 ? wdata[5:4] : PRV1; // @[CSR.scala 361:38 CSR.scala 362:14 CSR.scala 148:21]
  wire  _GEN_222 = csr_addr == 12'h300 ? wdata[3] : IE1; // @[CSR.scala 361:38 CSR.scala 363:14 CSR.scala 152:20]
  wire [1:0] _GEN_223 = csr_addr == 12'h300 ? wdata[2:1] : PRV; // @[CSR.scala 361:38 CSR.scala 364:14 CSR.scala 147:21]
  wire  _GEN_224 = csr_addr == 12'h300 ? wdata[0] : IE; // @[CSR.scala 361:38 CSR.scala 365:14 CSR.scala 151:20]
  wire  _GEN_225 = csr_addr == 12'h300 ? _GEN_6 : _GEN_201; // @[CSR.scala 361:38]
  wire  _GEN_226 = csr_addr == 12'h300 ? MSIP : _GEN_202; // @[CSR.scala 361:38 CSR.scala 174:21]
  wire  _GEN_227 = csr_addr == 12'h300 ? MTIE : _GEN_203; // @[CSR.scala 361:38 CSR.scala 171:21]
  wire  _GEN_228 = csr_addr == 12'h300 ? MSIE : _GEN_204; // @[CSR.scala 361:38 CSR.scala 177:21]
  wire [31:0] _GEN_229 = csr_addr == 12'h300 ? _GEN_4 : _GEN_205; // @[CSR.scala 361:38]
  wire [31:0] _GEN_230 = csr_addr == 12'h300 ? _GEN_5 : _GEN_206; // @[CSR.scala 361:38]
  wire [31:0] _GEN_231 = csr_addr == 12'h300 ? mtimecmp : _GEN_207; // @[CSR.scala 361:38 CSR.scala 185:21]
  wire [31:0] _GEN_232 = csr_addr == 12'h300 ? mscratch : _GEN_208; // @[CSR.scala 361:38 CSR.scala 187:21]
  wire [34:0] _GEN_233 = csr_addr == 12'h300 ? {{3'd0}, mepc} : _GEN_209; // @[CSR.scala 361:38 CSR.scala 189:17]
  wire [31:0] _GEN_234 = csr_addr == 12'h300 ? mcause : _GEN_210; // @[CSR.scala 361:38 CSR.scala 190:19]
  wire [31:0] _GEN_235 = csr_addr == 12'h300 ? mbadaddr : _GEN_211; // @[CSR.scala 361:38 CSR.scala 191:21]
  wire [31:0] _GEN_236 = csr_addr == 12'h300 ? mtohost : _GEN_212; // @[CSR.scala 361:38 CSR.scala 193:24]
  wire [31:0] _GEN_237 = csr_addr == 12'h300 ? mfromhost : _GEN_213; // @[CSR.scala 361:38]
  wire [31:0] _GEN_238 = csr_addr == 12'h300 ? _T_278 : _GEN_214; // @[CSR.scala 361:38 CSR.scala 320:9]
  wire [31:0] _GEN_239 = csr_addr == 12'h300 ? _GEN_8 : _GEN_215; // @[CSR.scala 361:38]
  wire [31:0] _GEN_240 = csr_addr == 12'h300 ? _GEN_7 : _GEN_216; // @[CSR.scala 361:38]
  wire [31:0] _GEN_241 = csr_addr == 12'h300 ? _GEN_9 : _GEN_217; // @[CSR.scala 361:38]
  wire [31:0] _GEN_242 = csr_addr == 12'h300 ? satp : _GEN_218; // @[CSR.scala 361:38 CSR.scala 202:21]
  wire [31:0] _GEN_243 = csr_addr == 12'h300 ? vmSwitchPC : _GEN_219; // @[CSR.scala 361:38 CSR.scala 289:27]
  wire [31:0] _GEN_244 = csr_addr == 12'h300 ? mtvec : _GEN_220; // @[CSR.scala 361:38 CSR.scala 164:24]
  wire [1:0] _GEN_245 = wen ? _GEN_221 : PRV1; // @[CSR.scala 360:21 CSR.scala 148:21]
  wire  _GEN_246 = wen ? _GEN_222 : IE1; // @[CSR.scala 360:21 CSR.scala 152:20]
  wire [1:0] _GEN_247 = wen ? _GEN_223 : PRV; // @[CSR.scala 360:21 CSR.scala 147:21]
  wire  _GEN_248 = wen ? _GEN_224 : IE; // @[CSR.scala 360:21 CSR.scala 151:20]
  wire  _GEN_249 = wen ? _GEN_225 : _GEN_6; // @[CSR.scala 360:21]
  wire  _GEN_250 = wen ? _GEN_226 : MSIP; // @[CSR.scala 360:21 CSR.scala 174:21]
  wire  _GEN_251 = wen ? _GEN_227 : MTIE; // @[CSR.scala 360:21 CSR.scala 171:21]
  wire  _GEN_252 = wen ? _GEN_228 : MSIE; // @[CSR.scala 360:21 CSR.scala 177:21]
  wire [31:0] _GEN_253 = wen ? _GEN_229 : _GEN_4; // @[CSR.scala 360:21]
  wire [31:0] _GEN_254 = wen ? _GEN_230 : _GEN_5; // @[CSR.scala 360:21]
  wire [34:0] _GEN_257 = wen ? _GEN_233 : {{3'd0}, mepc}; // @[CSR.scala 360:21 CSR.scala 189:17]
  wire [31:0] _GEN_260 = wen ? _GEN_236 : mtohost; // @[CSR.scala 360:21 CSR.scala 193:24]
  wire [31:0] _GEN_262 = wen ? _GEN_238 : _T_278; // @[CSR.scala 360:21 CSR.scala 320:9]
  wire [31:0] _GEN_263 = wen ? _GEN_239 : _GEN_8; // @[CSR.scala 360:21]
  wire [31:0] _GEN_264 = wen ? _GEN_240 : _GEN_7; // @[CSR.scala 360:21]
  wire [31:0] _GEN_265 = wen ? _GEN_241 : _GEN_9; // @[CSR.scala 360:21]
  wire [31:0] _GEN_266 = wen ? _GEN_242 : satp; // @[CSR.scala 360:21 CSR.scala 202:21]
  wire [31:0] _GEN_267 = wen ? _GEN_243 : vmSwitchPC; // @[CSR.scala 360:21 CSR.scala 289:27]
  wire [31:0] _GEN_268 = wen ? _GEN_244 : mtvec; // @[CSR.scala 360:21 CSR.scala 164:24]
  wire  _GEN_272 = isEret | _GEN_246; // @[CSR.scala 355:24 CSR.scala 359:12]
  wire [34:0] _GEN_281 = isEret ? {{3'd0}, mepc} : _GEN_257; // @[CSR.scala 355:24 CSR.scala 189:17]
  wire [34:0] _GEN_293 = io__expt ? {{3'd0}, _T_296} : _GEN_281; // @[CSR.scala 327:19 CSR.scala 328:14]
  wire  _GEN_301 = io__expt & _T_317; // @[CSR.scala 327:19]
  wire [34:0] _GEN_319 = _T_287 ? _GEN_293 : {{3'd0}, mepc}; // @[CSR.scala 326:19 CSR.scala 189:17]
  wire  clearPageFault = _T_287 & _GEN_301; // @[CSR.scala 326:19]
  assign io__out = _T_2 ? cycle : _T_92; // @[Lookup.scala 33:37]
  assign io__expt = t_expt | isDFCAct | writeDFCInvalid; // @[CSR.scala 309:34]
  assign io__evec = mtvec; // @[CSR.scala 311:11]
  assign io__epc = mepc; // @[CSR.scala 312:11]
  assign io__vmSwitch = csr_addr == 12'h180 & wen; // @[CSR.scala 288:40]
  assign io__vmSwitchPC = io__stall ? vmSwitchPC : io__pc; // @[CSR.scala 290:23]
  assign io__dfc_full = dfc_full_reg; // @[CSR.scala 226:15]
  assign io_vmSwitch = io__vmSwitch;
  assign io_in = io__in;
  assign clearPageFault_0 = clearPageFault;
  assign satp_0 = satp;
  always @(posedge clock) begin
    if (reset) begin // @[CSR.scala 132:25]
      time_ <= 32'h0; // @[CSR.scala 132:25]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (io__expt) begin // @[CSR.scala 327:19]
        time_ <= _GEN_4;
      end else if (isEret) begin // @[CSR.scala 355:24]
        time_ <= _GEN_4;
      end else begin
        time_ <= _GEN_253;
      end
    end else begin
      time_ <= _GEN_4;
    end
    if (reset) begin // @[CSR.scala 133:25]
      counter <= 32'h0; // @[CSR.scala 133:25]
    end else begin
      counter <= _T_268; // @[CSR.scala 315:11]
    end
    if (reset) begin // @[CSR.scala 134:25]
      timeh <= 32'h0; // @[CSR.scala 134:25]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (io__expt) begin // @[CSR.scala 327:19]
        timeh <= _GEN_5;
      end else if (isEret) begin // @[CSR.scala 355:24]
        timeh <= _GEN_5;
      end else begin
        timeh <= _GEN_254;
      end
    end else begin
      timeh <= _GEN_5;
    end
    if (reset) begin // @[CSR.scala 135:25]
      cycle <= 32'h0; // @[CSR.scala 135:25]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (io__expt) begin // @[CSR.scala 327:19]
        cycle <= _T_278; // @[CSR.scala 320:9]
      end else if (isEret) begin // @[CSR.scala 355:24]
        cycle <= _T_278; // @[CSR.scala 320:9]
      end else begin
        cycle <= _GEN_262;
      end
    end else begin
      cycle <= _T_278; // @[CSR.scala 320:9]
    end
    if (reset) begin // @[CSR.scala 136:25]
      cycleh <= 32'h0; // @[CSR.scala 136:25]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (io__expt) begin // @[CSR.scala 327:19]
        cycleh <= _GEN_7;
      end else if (isEret) begin // @[CSR.scala 355:24]
        cycleh <= _GEN_7;
      end else begin
        cycleh <= _GEN_264;
      end
    end else begin
      cycleh <= _GEN_7;
    end
    if (reset) begin // @[CSR.scala 137:25]
      instret <= 32'h0; // @[CSR.scala 137:25]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (io__expt) begin // @[CSR.scala 327:19]
        instret <= _GEN_8;
      end else if (isEret) begin // @[CSR.scala 355:24]
        instret <= _GEN_8;
      end else begin
        instret <= _GEN_263;
      end
    end else begin
      instret <= _GEN_8;
    end
    if (reset) begin // @[CSR.scala 138:25]
      instreth <= 32'h0; // @[CSR.scala 138:25]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (io__expt) begin // @[CSR.scala 327:19]
        instreth <= _GEN_9;
      end else if (isEret) begin // @[CSR.scala 355:24]
        instreth <= _GEN_9;
      end else begin
        instreth <= _GEN_265;
      end
    end else begin
      instreth <= _GEN_9;
    end
    if (reset) begin // @[CSR.scala 147:21]
      PRV <= 2'h3; // @[CSR.scala 147:21]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (io__expt) begin // @[CSR.scala 327:19]
        PRV <= 2'h3; // @[CSR.scala 347:12]
      end else if (isEret) begin // @[CSR.scala 355:24]
        PRV <= PRV1; // @[CSR.scala 356:12]
      end else begin
        PRV <= _GEN_247;
      end
    end
    if (reset) begin // @[CSR.scala 148:21]
      PRV1 <= 2'h3; // @[CSR.scala 148:21]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (io__expt) begin // @[CSR.scala 327:19]
        PRV1 <= PRV; // @[CSR.scala 349:12]
      end else if (isEret) begin // @[CSR.scala 355:24]
        PRV1 <= 2'h0; // @[CSR.scala 358:12]
      end else begin
        PRV1 <= _GEN_245;
      end
    end
    if (reset) begin // @[CSR.scala 151:20]
      IE <= 1'h0; // @[CSR.scala 151:20]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (io__expt) begin // @[CSR.scala 327:19]
        IE <= 1'h0; // @[CSR.scala 348:12]
      end else if (isEret) begin // @[CSR.scala 355:24]
        IE <= IE1; // @[CSR.scala 357:12]
      end else begin
        IE <= _GEN_248;
      end
    end
    if (reset) begin // @[CSR.scala 152:20]
      IE1 <= 1'h0; // @[CSR.scala 152:20]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (io__expt) begin // @[CSR.scala 327:19]
        IE1 <= IE; // @[CSR.scala 350:12]
      end else begin
        IE1 <= _GEN_272;
      end
    end
    if (reset) begin // @[CSR.scala 164:24]
      mtvec <= 32'h100; // @[CSR.scala 164:24]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (!(io__expt)) begin // @[CSR.scala 327:19]
        if (!(isEret)) begin // @[CSR.scala 355:24]
          mtvec <= _GEN_268;
        end
      end
    end
    if (reset) begin // @[CSR.scala 168:21]
      MTIP <= 1'h0; // @[CSR.scala 168:21]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (io__expt) begin // @[CSR.scala 327:19]
        MTIP <= _GEN_6;
      end else if (isEret) begin // @[CSR.scala 355:24]
        MTIP <= _GEN_6;
      end else begin
        MTIP <= _GEN_249;
      end
    end else begin
      MTIP <= _GEN_6;
    end
    if (reset) begin // @[CSR.scala 171:21]
      MTIE <= 1'h0; // @[CSR.scala 171:21]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (!(io__expt)) begin // @[CSR.scala 327:19]
        if (!(isEret)) begin // @[CSR.scala 355:24]
          MTIE <= _GEN_251;
        end
      end
    end
    if (reset) begin // @[CSR.scala 174:21]
      MSIP <= 1'h0; // @[CSR.scala 174:21]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (!(io__expt)) begin // @[CSR.scala 327:19]
        if (!(isEret)) begin // @[CSR.scala 355:24]
          MSIP <= _GEN_250;
        end
      end
    end
    if (reset) begin // @[CSR.scala 177:21]
      MSIE <= 1'h0; // @[CSR.scala 177:21]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (!(io__expt)) begin // @[CSR.scala 327:19]
        if (!(isEret)) begin // @[CSR.scala 355:24]
          MSIE <= _GEN_252;
        end
      end
    end
    if (reset) begin // @[CSR.scala 183:37]
      uartInterruptPending <= 1'h0; // @[CSR.scala 183:37]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (io__expt) begin // @[CSR.scala 327:19]
        if (isUartInterrupt) begin // @[CSR.scala 353:28]
          uartInterruptPending <= 1'h0; // @[CSR.scala 353:50]
        end else begin
          uartInterruptPending <= _GEN_1;
        end
      end else begin
        uartInterruptPending <= _GEN_1;
      end
    end else begin
      uartInterruptPending <= _GEN_1;
    end
    if (_T_287) begin // @[CSR.scala 326:19]
      if (!(io__expt)) begin // @[CSR.scala 327:19]
        if (!(isEret)) begin // @[CSR.scala 355:24]
          if (wen) begin // @[CSR.scala 360:21]
            mtimecmp <= _GEN_231;
          end
        end
      end
    end
    if (_T_287) begin // @[CSR.scala 326:19]
      if (!(io__expt)) begin // @[CSR.scala 327:19]
        if (!(isEret)) begin // @[CSR.scala 355:24]
          if (wen) begin // @[CSR.scala 360:21]
            mscratch <= _GEN_232;
          end
        end
      end
    end
    mepc <= _GEN_319[31:0];
    if (_T_287) begin // @[CSR.scala 326:19]
      if (io__expt) begin // @[CSR.scala 327:19]
        if (isDFCAct) begin // @[CSR.scala 331:20]
          mcause <= 32'h12;
        end else if (iaddrInvalid) begin // @[CSR.scala 332:20]
          mcause <= 32'h0;
        end else begin
          mcause <= _T_308;
        end
      end else if (!(isEret)) begin // @[CSR.scala 355:24]
        if (wen) begin // @[CSR.scala 360:21]
          mcause <= _GEN_234;
        end
      end
    end
    if (_T_287) begin // @[CSR.scala 326:19]
      if (io__expt) begin // @[CSR.scala 327:19]
        if (iaddrInvalid | laddrInvalid | saddrInvalid | isInstructionFault | isLoadFault | isStoreFault) begin // @[CSR.scala 352:111]
          mbadaddr <= io__addr; // @[CSR.scala 352:122]
        end
      end else if (!(isEret)) begin // @[CSR.scala 355:24]
        if (wen) begin // @[CSR.scala 360:21]
          mbadaddr <= _GEN_235;
        end
      end
    end
    if (reset) begin // @[CSR.scala 193:24]
      mtohost <= 32'h0; // @[CSR.scala 193:24]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (!(io__expt)) begin // @[CSR.scala 327:19]
        if (!(isEret)) begin // @[CSR.scala 355:24]
          mtohost <= _GEN_260;
        end
      end
    end
    if (_T_287) begin // @[CSR.scala 326:19]
      if (!(io__expt)) begin // @[CSR.scala 327:19]
        if (!(isEret)) begin // @[CSR.scala 355:24]
          if (wen) begin // @[CSR.scala 360:21]
            mfromhost <= _GEN_237;
          end
        end
      end
    end
    if (reset) begin // @[CSR.scala 202:21]
      satp <= 32'h0; // @[CSR.scala 202:21]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (!(io__expt)) begin // @[CSR.scala 327:19]
        if (!(isEret)) begin // @[CSR.scala 355:24]
          satp <= _GEN_266;
        end
      end
    end
    if (reset) begin // @[CSR.scala 224:24]
      dfc_pid <= 32'h0; // @[CSR.scala 224:24]
    end else if (isDFCAct) begin // @[CSR.scala 299:17]
      dfc_pid <= {{16'd0}, io__dfc_pid}; // @[CSR.scala 300:13]
    end
    if (reset) begin // @[CSR.scala 225:29]
      dfc_full_reg <= 1'h0; // @[CSR.scala 225:29]
    end else if (io__table_f_data_valid) begin // @[CSR.scala 302:30]
      dfc_full_reg <= io__table_f_data_bits_full_sig; // @[CSR.scala 303:18]
    end
    if (reset) begin // @[CSR.scala 289:27]
      vmSwitchPC <= 32'h0; // @[CSR.scala 289:27]
    end else if (_T_287) begin // @[CSR.scala 326:19]
      if (!(io__expt)) begin // @[CSR.scala 327:19]
        if (!(isEret)) begin // @[CSR.scala 355:24]
          vmSwitchPC <= _GEN_267;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  time_ = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  timeh = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  cycle = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  cycleh = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  instret = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  instreth = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  PRV = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  PRV1 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  IE = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  IE1 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  mtvec = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  MTIP = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  MTIE = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  MSIP = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  MSIE = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  uartInterruptPending = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  mtimecmp = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  mscratch = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  mepc = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  mcause = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  mbadaddr = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  mtohost = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  mfromhost = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  satp = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  dfc_pid = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  dfc_full_reg = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  vmSwitchPC = _RAND_27[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegFile(
  input         clock,
  input  [4:0]  io_raddr1,
  input  [4:0]  io_raddr2,
  output [31:0] io_rdata1,
  output [31:0] io_rdata2,
  input         io_wen,
  input  [4:0]  io_waddr,
  input  [31:0] io_wdata
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [31:0] regs [0:31]; // @[RegFile.scala 25:17]
  wire [31:0] regs_MPORT_data; // @[RegFile.scala 25:17]
  wire [4:0] regs_MPORT_addr; // @[RegFile.scala 25:17]
  wire [31:0] regs_MPORT_1_data; // @[RegFile.scala 25:17]
  wire [4:0] regs_MPORT_1_addr; // @[RegFile.scala 25:17]
  wire [31:0] regs_MPORT_2_data; // @[RegFile.scala 25:17]
  wire [4:0] regs_MPORT_2_addr; // @[RegFile.scala 25:17]
  wire  regs_MPORT_2_mask; // @[RegFile.scala 25:17]
  wire  regs_MPORT_2_en; // @[RegFile.scala 25:17]
  wire  _T_4 = |io_waddr; // @[RegFile.scala 29:26]
  assign regs_MPORT_addr = io_raddr1;
  assign regs_MPORT_data = regs[regs_MPORT_addr]; // @[RegFile.scala 25:17]
  assign regs_MPORT_1_addr = io_raddr2;
  assign regs_MPORT_1_data = regs[regs_MPORT_1_addr]; // @[RegFile.scala 25:17]
  assign regs_MPORT_2_data = io_wdata;
  assign regs_MPORT_2_addr = io_waddr;
  assign regs_MPORT_2_mask = 1'h1;
  assign regs_MPORT_2_en = io_wen & _T_4;
  assign io_rdata1 = |io_raddr1 ? regs_MPORT_data : 32'h0; // @[RegFile.scala 27:19]
  assign io_rdata2 = |io_raddr2 ? regs_MPORT_1_data : 32'h0; // @[RegFile.scala 28:19]
  always @(posedge clock) begin
    if(regs_MPORT_2_en & regs_MPORT_2_mask) begin
      regs[regs_MPORT_2_addr] <= regs_MPORT_2_data; // @[RegFile.scala 25:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regs[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ALUArea(
  input  [31:0] io_A,
  input  [31:0] io_B,
  input  [3:0]  io_alu_op,
  output [31:0] io_out,
  output [31:0] io_sum
);
  wire [31:0] _T_2 = 32'h0 - io_B; // @[ALU.scala 63:38]
  wire [31:0] _T_3 = io_alu_op[0] ? _T_2 : io_B; // @[ALU.scala 63:23]
  wire [31:0] sum = io_A + _T_3; // @[ALU.scala 63:18]
  wire  _T_12 = io_alu_op[1] ? io_B[31] : io_A[31]; // @[ALU.scala 65:16]
  wire  cmp = io_A[31] == io_B[31] ? sum[31] : _T_12; // @[ALU.scala 64:16]
  wire [4:0] shamt = io_B[4:0]; // @[ALU.scala 66:20]
  wire [31:0] _T_17 = {{16'd0}, io_A[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_19 = {io_A[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_21 = _T_19 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_22 = _T_17 | _T_21; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_0 = {{8'd0}, _T_22[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_27 = _GEN_0 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_29 = {_T_22[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_31 = _T_29 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_32 = _T_27 | _T_31; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_1 = {{4'd0}, _T_32[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_37 = _GEN_1 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_39 = {_T_32[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_41 = _T_39 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_42 = _T_37 | _T_41; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_2 = {{2'd0}, _T_42[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_47 = _GEN_2 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_49 = {_T_42[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_51 = _T_49 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_52 = _T_47 | _T_51; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_3 = {{1'd0}, _T_52[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_57 = _GEN_3 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_59 = {_T_52[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_61 = _T_59 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] _T_62 = _T_57 | _T_61; // @[Bitwise.scala 103:39]
  wire [31:0] shin = io_alu_op[3] ? io_A : _T_62; // @[ALU.scala 67:19]
  wire  hi = io_alu_op[0] & shin[31]; // @[ALU.scala 68:34]
  wire [32:0] _T_66 = {hi,shin}; // @[ALU.scala 68:57]
  wire [32:0] _T_67 = $signed(_T_66) >>> shamt; // @[ALU.scala 68:64]
  wire [31:0] shiftr = _T_67[31:0]; // @[ALU.scala 68:73]
  wire [31:0] _T_71 = {{16'd0}, shiftr[31:16]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_73 = {shiftr[15:0], 16'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_75 = _T_73 & 32'hffff0000; // @[Bitwise.scala 103:75]
  wire [31:0] _T_76 = _T_71 | _T_75; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_4 = {{8'd0}, _T_76[31:8]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_81 = _GEN_4 & 32'hff00ff; // @[Bitwise.scala 103:31]
  wire [31:0] _T_83 = {_T_76[23:0], 8'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_85 = _T_83 & 32'hff00ff00; // @[Bitwise.scala 103:75]
  wire [31:0] _T_86 = _T_81 | _T_85; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_5 = {{4'd0}, _T_86[31:4]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_91 = _GEN_5 & 32'hf0f0f0f; // @[Bitwise.scala 103:31]
  wire [31:0] _T_93 = {_T_86[27:0], 4'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_95 = _T_93 & 32'hf0f0f0f0; // @[Bitwise.scala 103:75]
  wire [31:0] _T_96 = _T_91 | _T_95; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_6 = {{2'd0}, _T_96[31:2]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_101 = _GEN_6 & 32'h33333333; // @[Bitwise.scala 103:31]
  wire [31:0] _T_103 = {_T_96[29:0], 2'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_105 = _T_103 & 32'hcccccccc; // @[Bitwise.scala 103:75]
  wire [31:0] _T_106 = _T_101 | _T_105; // @[Bitwise.scala 103:39]
  wire [31:0] _GEN_7 = {{1'd0}, _T_106[31:1]}; // @[Bitwise.scala 103:31]
  wire [31:0] _T_111 = _GEN_7 & 32'h55555555; // @[Bitwise.scala 103:31]
  wire [31:0] _T_113 = {_T_106[30:0], 1'h0}; // @[Bitwise.scala 103:65]
  wire [31:0] _T_115 = _T_113 & 32'haaaaaaaa; // @[Bitwise.scala 103:75]
  wire [31:0] shiftl = _T_111 | _T_115; // @[Bitwise.scala 103:39]
  wire [31:0] _T_127 = io_A & io_B; // @[ALU.scala 76:38]
  wire [31:0] _T_129 = io_A | io_B; // @[ALU.scala 77:38]
  wire [31:0] _T_131 = io_A ^ io_B; // @[ALU.scala 78:38]
  wire [31:0] _T_133 = io_alu_op == 4'ha ? io_A : io_B; // @[ALU.scala 79:8]
  wire [31:0] _T_134 = io_alu_op == 4'h4 ? _T_131 : _T_133; // @[ALU.scala 78:8]
  wire [31:0] _T_135 = io_alu_op == 4'h3 ? _T_129 : _T_134; // @[ALU.scala 77:8]
  wire [31:0] _T_136 = io_alu_op == 4'h2 ? _T_127 : _T_135; // @[ALU.scala 76:8]
  wire [31:0] _T_137 = io_alu_op == 4'h6 ? shiftl : _T_136; // @[ALU.scala 75:8]
  wire [31:0] _T_138 = io_alu_op == 4'h9 | io_alu_op == 4'h8 ? shiftr : _T_137; // @[ALU.scala 74:8]
  wire [31:0] _T_139 = io_alu_op == 4'h5 | io_alu_op == 4'h7 ? {{31'd0}, cmp} : _T_138; // @[ALU.scala 73:8]
  assign io_out = io_alu_op == 4'h0 | io_alu_op == 4'h1 ? sum : _T_139; // @[ALU.scala 72:8]
  assign io_sum = io_A + _T_3; // @[ALU.scala 63:18]
endmodule
module ImmGenWire(
  input  [31:0] io_inst,
  input  [2:0]  io_sel,
  output [31:0] io_out
);
  wire [11:0] Iimm = io_inst[31:20]; // @[ImmGen.scala 28:30]
  wire [6:0] hi = io_inst[31:25]; // @[ImmGen.scala 29:25]
  wire [4:0] lo = io_inst[11:7]; // @[ImmGen.scala 29:42]
  wire [11:0] Simm = {hi,lo}; // @[ImmGen.scala 29:50]
  wire  hi_hi_hi = io_inst[31]; // @[ImmGen.scala 30:25]
  wire  hi_hi_lo = io_inst[7]; // @[ImmGen.scala 30:38]
  wire [5:0] hi_lo = io_inst[30:25]; // @[ImmGen.scala 30:50]
  wire [3:0] lo_hi = io_inst[11:8]; // @[ImmGen.scala 30:67]
  wire [12:0] Bimm = {hi_hi_hi,hi_hi_lo,hi_lo,lo_hi,1'h0}; // @[ImmGen.scala 30:86]
  wire [19:0] hi_2 = io_inst[31:12]; // @[ImmGen.scala 31:25]
  wire [31:0] Uimm = {hi_2,12'h0}; // @[ImmGen.scala 31:46]
  wire [7:0] hi_hi_lo_1 = io_inst[19:12]; // @[ImmGen.scala 32:38]
  wire  hi_lo_1 = io_inst[20]; // @[ImmGen.scala 32:55]
  wire [3:0] lo_hi_lo = io_inst[24:21]; // @[ImmGen.scala 32:85]
  wire [20:0] Jimm = {hi_hi_hi,hi_hi_lo_1,hi_lo_1,hi_lo,lo_hi_lo,1'h0}; // @[ImmGen.scala 32:105]
  wire [5:0] Zimm = {1'b0,$signed(io_inst[19:15])}; // @[ImmGen.scala 33:30]
  wire [11:0] _T_7 = $signed(Iimm) & -12'sh2; // @[ImmGen.scala 35:36]
  wire [11:0] _T_9 = 3'h1 == io_sel ? $signed(Iimm) : $signed(_T_7); // @[Mux.scala 80:57]
  wire [11:0] _T_11 = 3'h2 == io_sel ? $signed(Simm) : $signed(_T_9); // @[Mux.scala 80:57]
  wire [12:0] _T_13 = 3'h5 == io_sel ? $signed(Bimm) : $signed({{1{_T_11[11]}},_T_11}); // @[Mux.scala 80:57]
  wire [31:0] _T_15 = 3'h3 == io_sel ? $signed(Uimm) : $signed({{19{_T_13[12]}},_T_13}); // @[Mux.scala 80:57]
  wire [31:0] _T_17 = 3'h4 == io_sel ? $signed({{11{Jimm[20]}},Jimm}) : $signed(_T_15); // @[Mux.scala 80:57]
  assign io_out = 3'h6 == io_sel ? $signed({{26{Zimm[5]}},Zimm}) : $signed(_T_17); // @[ImmGen.scala 36:100]
endmodule
module BrCondArea(
  input  [31:0] io_rs1,
  input  [31:0] io_rs2,
  input  [2:0]  io_br_type,
  output        io_taken
);
  wire [31:0] diff = io_rs1 - io_rs2; // @[BrCond.scala 44:21]
  wire  neq = |diff; // @[BrCond.scala 45:19]
  wire  eq = ~neq; // @[BrCond.scala 46:14]
  wire  isSameSign = io_rs1[31] == io_rs2[31]; // @[BrCond.scala 47:35]
  wire  lt = isSameSign ? diff[31] : io_rs1[31]; // @[BrCond.scala 48:17]
  wire  ltu = isSameSign ? diff[31] : io_rs2[31]; // @[BrCond.scala 49:17]
  wire  ge = ~lt; // @[BrCond.scala 50:14]
  wire  geu = ~ltu; // @[BrCond.scala 51:14]
  wire  _T_10 = io_br_type == 3'h6 & neq; // @[BrCond.scala 54:29]
  wire  _T_11 = io_br_type == 3'h3 & eq | _T_10; // @[BrCond.scala 53:36]
  wire  _T_13 = io_br_type == 3'h2 & lt; // @[BrCond.scala 55:29]
  wire  _T_14 = _T_11 | _T_13; // @[BrCond.scala 54:37]
  wire  _T_16 = io_br_type == 3'h5 & ge; // @[BrCond.scala 56:29]
  wire  _T_17 = _T_14 | _T_16; // @[BrCond.scala 55:36]
  wire  _T_19 = io_br_type == 3'h1 & ltu; // @[BrCond.scala 57:30]
  wire  _T_20 = _T_17 | _T_19; // @[BrCond.scala 56:36]
  wire  _T_22 = io_br_type == 3'h4 & geu; // @[BrCond.scala 58:30]
  assign io_taken = _T_20 | _T_22; // @[BrCond.scala 57:38]
endmodule
module Datapath(
  input         clock,
  input         reset,
  output        io_icache_req_valid,
  output [31:0] io_icache_req_bits_addr,
  input         io_icache_resp_valid,
  input  [31:0] io_icache_resp_bits_data,
  output        io_dcache_abort,
  output        io_dcache_req_valid,
  output [31:0] io_dcache_req_bits_addr,
  output [31:0] io_dcache_req_bits_data,
  output [3:0]  io_dcache_req_bits_mask,
  input         io_dcache_resp_valid,
  input  [31:0] io_dcache_resp_bits_data,
  output [31:0] io_ctrl_inst,
  input  [1:0]  io_ctrl_pc_sel,
  input         io_ctrl_inst_kill,
  input         io_ctrl_A_sel,
  input         io_ctrl_B_sel,
  input  [2:0]  io_ctrl_imm_sel,
  input  [3:0]  io_ctrl_alu_op,
  input  [2:0]  io_ctrl_br_type,
  input  [1:0]  io_ctrl_st_type,
  input  [2:0]  io_ctrl_ld_type,
  input  [1:0]  io_ctrl_wb_sel,
  input         io_ctrl_wb_en,
  input  [2:0]  io_ctrl_csr_cmd,
  input         io_ctrl_illegal,
  input  [2:0]  io_ctrl_dfc_cmd,
  output        io_table_w_data_valid,
  output [31:0] io_table_w_data_bits_listenAddr,
  output [15:0] io_table_w_data_bits_wPid,
  output        io_table_l_data_valid,
  output [31:0] io_table_l_data_bits_listenAddr,
  output        io_table_e_data_ready,
  input         io_table_e_data_valid,
  input  [15:0] io_table_e_data_bits_pid,
  input         io_table_f_data_valid,
  input         io_table_f_data_bits_full_sig,
  input         io_rxChannel_valid,
  input  [1:0]  pageFault,
  output        io_vmSwitch,
  output [31:0] io_in,
  output        clearPageFault,
  input  [1:0]  pageFault_0,
  output [31:0] satp
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  csr_clock; // @[Datapath.scala 29:23]
  wire  csr_reset; // @[Datapath.scala 29:23]
  wire  csr_io__stall; // @[Datapath.scala 29:23]
  wire [2:0] csr_io__cmd; // @[Datapath.scala 29:23]
  wire [31:0] csr_io__in; // @[Datapath.scala 29:23]
  wire [31:0] csr_io__out; // @[Datapath.scala 29:23]
  wire [31:0] csr_io__pc; // @[Datapath.scala 29:23]
  wire [31:0] csr_io__addr; // @[Datapath.scala 29:23]
  wire [31:0] csr_io__inst; // @[Datapath.scala 29:23]
  wire  csr_io__illegal; // @[Datapath.scala 29:23]
  wire [1:0] csr_io__st_type; // @[Datapath.scala 29:23]
  wire [2:0] csr_io__ld_type; // @[Datapath.scala 29:23]
  wire  csr_io__pc_check; // @[Datapath.scala 29:23]
  wire  csr_io__expt; // @[Datapath.scala 29:23]
  wire [31:0] csr_io__evec; // @[Datapath.scala 29:23]
  wire [31:0] csr_io__epc; // @[Datapath.scala 29:23]
  wire  csr_io__vmSwitch; // @[Datapath.scala 29:23]
  wire [31:0] csr_io__vmSwitchPC; // @[Datapath.scala 29:23]
  wire [2:0] csr_io__dfc_cmd; // @[Datapath.scala 29:23]
  wire [15:0] csr_io__dfc_pid; // @[Datapath.scala 29:23]
  wire  csr_io__table_f_data_valid; // @[Datapath.scala 29:23]
  wire  csr_io__table_f_data_bits_full_sig; // @[Datapath.scala 29:23]
  wire  csr_io__dfc_full; // @[Datapath.scala 29:23]
  wire  csr_uartRxValid_0; // @[Datapath.scala 29:23]
  wire [1:0] csr_dmmu; // @[Datapath.scala 29:23]
  wire  csr_io_vmSwitch; // @[Datapath.scala 29:23]
  wire [31:0] csr_io_in; // @[Datapath.scala 29:23]
  wire  csr_clearPageFault_0; // @[Datapath.scala 29:23]
  wire [1:0] csr_immu; // @[Datapath.scala 29:23]
  wire [31:0] csr_satp_0; // @[Datapath.scala 29:23]
  wire  regFile_clock; // @[Datapath.scala 30:23]
  wire [4:0] regFile_io_raddr1; // @[Datapath.scala 30:23]
  wire [4:0] regFile_io_raddr2; // @[Datapath.scala 30:23]
  wire [31:0] regFile_io_rdata1; // @[Datapath.scala 30:23]
  wire [31:0] regFile_io_rdata2; // @[Datapath.scala 30:23]
  wire  regFile_io_wen; // @[Datapath.scala 30:23]
  wire [4:0] regFile_io_waddr; // @[Datapath.scala 30:23]
  wire [31:0] regFile_io_wdata; // @[Datapath.scala 30:23]
  wire [31:0] alu_io_A; // @[Config.scala 13:50]
  wire [31:0] alu_io_B; // @[Config.scala 13:50]
  wire [3:0] alu_io_alu_op; // @[Config.scala 13:50]
  wire [31:0] alu_io_out; // @[Config.scala 13:50]
  wire [31:0] alu_io_sum; // @[Config.scala 13:50]
  wire [31:0] immGen_io_inst; // @[Config.scala 14:50]
  wire [2:0] immGen_io_sel; // @[Config.scala 14:50]
  wire [31:0] immGen_io_out; // @[Config.scala 14:50]
  wire [31:0] brCond_io_rs1; // @[Config.scala 15:50]
  wire [31:0] brCond_io_rs2; // @[Config.scala 15:50]
  wire [2:0] brCond_io_br_type; // @[Config.scala 15:50]
  wire  brCond_io_taken; // @[Config.scala 15:50]
  reg [31:0] fe_inst; // @[Datapath.scala 40:24]
  reg [32:0] fe_pc; // @[Datapath.scala 41:20]
  reg [31:0] ew_inst; // @[Datapath.scala 44:24]
  reg [32:0] ew_pc; // @[Datapath.scala 45:20]
  reg [31:0] ew_alu; // @[Datapath.scala 46:20]
  reg [31:0] csr_in; // @[Datapath.scala 47:20]
  reg [1:0] st_type; // @[Datapath.scala 50:21]
  reg [2:0] ld_type; // @[Datapath.scala 51:21]
  reg [1:0] wb_sel; // @[Datapath.scala 52:21]
  reg  wb_en; // @[Datapath.scala 53:21]
  reg [2:0] csr_cmd; // @[Datapath.scala 54:21]
  reg  illegal; // @[Datapath.scala 55:21]
  reg  pc_check; // @[Datapath.scala 56:21]
  reg [2:0] csr_dfc_cmd; // @[Datapath.scala 59:24]
  reg  started; // @[Datapath.scala 62:24]
  wire  stall = ~io_icache_resp_valid | ~io_dcache_resp_valid; // @[Datapath.scala 63:37]
  wire [31:0] _T_4 = 32'h200 - 32'h4; // @[Datapath.scala 64:41]
  reg [32:0] pc; // @[Datapath.scala 64:21]
  wire  _T_6 = io_ctrl_pc_sel == 2'h1; // @[Datapath.scala 69:33]
  wire [31:0] _T_8 = {{1'd0}, alu_io_sum[31:1]}; // @[Datapath.scala 69:75]
  wire [32:0] _T_9 = {_T_8, 1'h0}; // @[Datapath.scala 69:82]
  wire [31:0] _T_12 = csr_io__vmSwitchPC + 32'h4; // @[Datapath.scala 71:52]
  wire [32:0] _T_14 = pc + 33'h4; // @[Datapath.scala 71:61]
  wire [32:0] _T_15 = csr_io__vmSwitch ? {{1'd0}, _T_12} : _T_14; // @[Datapath.scala 71:17]
  wire [32:0] _T_16 = io_ctrl_pc_sel == 2'h2 ? pc : _T_15; // @[Datapath.scala 70:17]
  wire [32:0] _T_17 = io_ctrl_pc_sel == 2'h1 | brCond_io_taken ? _T_9 : _T_16; // @[Datapath.scala 69:17]
  wire [32:0] _T_18 = io_ctrl_pc_sel == 2'h3 ? {{1'd0}, csr_io__epc} : _T_17; // @[Datapath.scala 68:17]
  wire [32:0] _T_19 = csr_io__expt ? {{1'd0}, csr_io__evec} : _T_18; // @[Datapath.scala 66:32]
  wire [32:0] npc = stall ? pc : _T_19; // @[Datapath.scala 66:17]
  wire  _T_24 = ~stall; // @[Datapath.scala 83:30]
  wire [4:0] rs1_addr = fe_inst[19:15]; // @[Datapath.scala 98:25]
  wire [4:0] rs2_addr = fe_inst[24:20]; // @[Datapath.scala 99:25]
  wire [4:0] wb_rd_addr = ew_inst[11:7]; // @[Datapath.scala 108:27]
  wire  rs1hazard = wb_en & |rs1_addr & rs1_addr == wb_rd_addr; // @[Datapath.scala 109:41]
  wire  rs2hazard = wb_en & |rs2_addr & rs2_addr == wb_rd_addr; // @[Datapath.scala 110:41]
  wire  _T_32 = wb_sel == 2'h0; // @[Datapath.scala 111:24]
  wire [31:0] rs1 = wb_sel == 2'h0 & rs1hazard ? ew_alu : regFile_io_rdata1; // @[Datapath.scala 111:16]
  wire [31:0] rs2 = _T_32 & rs2hazard ? ew_alu : regFile_io_rdata2; // @[Datapath.scala 112:16]
  wire [32:0] _T_37 = io_ctrl_A_sel ? {{1'd0}, rs1} : fe_pc; // @[Datapath.scala 115:18]
  wire [31:0] _T_40 = stall ? ew_alu : alu_io_sum; // @[Datapath.scala 125:20]
  wire [31:0] _T_41 = {{2'd0}, _T_40[31:2]}; // @[Datapath.scala 125:48]
  wire [33:0] _GEN_28 = {_T_41, 2'h0}; // @[Datapath.scala 125:55]
  wire [34:0] daddr = {{1'd0}, _GEN_28}; // @[Datapath.scala 125:55]
  wire [4:0] _GEN_29 = {alu_io_sum[1], 4'h0}; // @[Datapath.scala 126:31]
  wire [7:0] _T_43 = {{3'd0}, _GEN_29}; // @[Datapath.scala 126:31]
  wire [3:0] _T_45 = {alu_io_sum[0], 3'h0}; // @[Datapath.scala 126:54]
  wire [7:0] _GEN_30 = {{4'd0}, _T_45}; // @[Datapath.scala 126:38]
  wire [7:0] woffset = _T_43 | _GEN_30; // @[Datapath.scala 126:38]
  wire [286:0] _GEN_31 = {{255'd0}, rs2}; // @[Datapath.scala 129:34]
  wire [286:0] _T_51 = _GEN_31 << woffset; // @[Datapath.scala 129:34]
  wire [1:0] _T_52 = stall ? st_type : io_ctrl_st_type; // @[Datapath.scala 130:43]
  wire [4:0] _T_54 = 5'h3 << alu_io_sum[1:0]; // @[Datapath.scala 133:23]
  wire [3:0] _T_56 = 4'h1 << alu_io_sum[1:0]; // @[Datapath.scala 134:23]
  wire [3:0] _T_58 = 2'h1 == _T_52 ? 4'hf : 4'h0; // @[Mux.scala 80:57]
  wire [4:0] _T_60 = 2'h2 == _T_52 ? _T_54 : {{1'd0}, _T_58}; // @[Mux.scala 80:57]
  wire [4:0] _T_62 = 2'h3 == _T_52 ? {{1'd0}, _T_56} : _T_60; // @[Mux.scala 80:57]
  wire  _T_71 = ~csr_io__expt; // @[Datapath.scala 147:24]
  wire  _T_73 = ~csr_io__vmSwitch; // @[Datapath.scala 147:40]
  wire [4:0] _GEN_32 = {ew_alu[1], 4'h0}; // @[Datapath.scala 164:27]
  wire [7:0] _T_79 = {{3'd0}, _GEN_32}; // @[Datapath.scala 164:27]
  wire [3:0] _T_81 = {ew_alu[0], 3'h0}; // @[Datapath.scala 164:46]
  wire [7:0] _GEN_33 = {{4'd0}, _T_81}; // @[Datapath.scala 164:34]
  wire [7:0] loffset = _T_79 | _GEN_33; // @[Datapath.scala 164:34]
  wire [31:0] lshift = io_dcache_resp_bits_data >> loffset; // @[Datapath.scala 165:42]
  wire [32:0] _T_82 = {1'b0,$signed(io_dcache_resp_bits_data)}; // @[Datapath.scala 166:61]
  wire [15:0] _T_84 = lshift[15:0]; // @[Datapath.scala 167:29]
  wire [7:0] _T_86 = lshift[7:0]; // @[Datapath.scala 167:60]
  wire [16:0] _T_88 = {1'b0,$signed(lshift[15:0])}; // @[Datapath.scala 168:29]
  wire [8:0] _T_90 = {1'b0,$signed(lshift[7:0])}; // @[Datapath.scala 168:60]
  wire [32:0] _T_92 = 3'h2 == ld_type ? $signed({{17{_T_84[15]}},_T_84}) : $signed(_T_82); // @[Mux.scala 80:57]
  wire [32:0] _T_94 = 3'h3 == ld_type ? $signed({{25{_T_86[7]}},_T_86}) : $signed(_T_92); // @[Mux.scala 80:57]
  wire [32:0] _T_96 = 3'h4 == ld_type ? $signed({{16{_T_88[16]}},_T_88}) : $signed(_T_94); // @[Mux.scala 80:57]
  wire [32:0] load = 3'h5 == ld_type ? $signed({{24{_T_90[8]}},_T_90}) : $signed(_T_96); // @[Mux.scala 80:57]
  wire [32:0] _T_100 = {1'b0,$signed(ew_alu)}; // @[Datapath.scala 190:43]
  wire [32:0] _T_102 = ew_pc + 33'h4; // @[Datapath.scala 192:22]
  wire [33:0] _T_103 = {1'b0,$signed(_T_102)}; // @[Datapath.scala 192:29]
  wire [32:0] _T_104 = {1'b0,$signed(csr_io__out)}; // @[Datapath.scala 193:26]
  wire [32:0] _T_106 = 2'h1 == wb_sel ? $signed(load) : $signed(_T_100); // @[Mux.scala 80:57]
  wire [33:0] _T_108 = 2'h2 == wb_sel ? $signed(_T_103) : $signed({{1{_T_106[32]}},_T_106}); // @[Mux.scala 80:57]
  wire [33:0] regWrite = 2'h3 == wb_sel ? $signed({{1{_T_104[32]}},_T_104}) : $signed(_T_108); // @[Datapath.scala 193:34]
  CSR csr ( // @[Datapath.scala 29:23]
    .clock(csr_clock),
    .reset(csr_reset),
    .io__stall(csr_io__stall),
    .io__cmd(csr_io__cmd),
    .io__in(csr_io__in),
    .io__out(csr_io__out),
    .io__pc(csr_io__pc),
    .io__addr(csr_io__addr),
    .io__inst(csr_io__inst),
    .io__illegal(csr_io__illegal),
    .io__st_type(csr_io__st_type),
    .io__ld_type(csr_io__ld_type),
    .io__pc_check(csr_io__pc_check),
    .io__expt(csr_io__expt),
    .io__evec(csr_io__evec),
    .io__epc(csr_io__epc),
    .io__vmSwitch(csr_io__vmSwitch),
    .io__vmSwitchPC(csr_io__vmSwitchPC),
    .io__dfc_cmd(csr_io__dfc_cmd),
    .io__dfc_pid(csr_io__dfc_pid),
    .io__table_f_data_valid(csr_io__table_f_data_valid),
    .io__table_f_data_bits_full_sig(csr_io__table_f_data_bits_full_sig),
    .io__dfc_full(csr_io__dfc_full),
    .uartRxValid_0(csr_uartRxValid_0),
    .dmmu(csr_dmmu),
    .io_vmSwitch(csr_io_vmSwitch),
    .io_in(csr_io_in),
    .clearPageFault_0(csr_clearPageFault_0),
    .immu(csr_immu),
    .satp_0(csr_satp_0)
  );
  RegFile regFile ( // @[Datapath.scala 30:23]
    .clock(regFile_clock),
    .io_raddr1(regFile_io_raddr1),
    .io_raddr2(regFile_io_raddr2),
    .io_rdata1(regFile_io_rdata1),
    .io_rdata2(regFile_io_rdata2),
    .io_wen(regFile_io_wen),
    .io_waddr(regFile_io_waddr),
    .io_wdata(regFile_io_wdata)
  );
  ALUArea alu ( // @[Config.scala 13:50]
    .io_A(alu_io_A),
    .io_B(alu_io_B),
    .io_alu_op(alu_io_alu_op),
    .io_out(alu_io_out),
    .io_sum(alu_io_sum)
  );
  ImmGenWire immGen ( // @[Config.scala 14:50]
    .io_inst(immGen_io_inst),
    .io_sel(immGen_io_sel),
    .io_out(immGen_io_out)
  );
  BrCondArea brCond ( // @[Config.scala 15:50]
    .io_rs1(brCond_io_rs1),
    .io_rs2(brCond_io_rs2),
    .io_br_type(brCond_io_br_type),
    .io_taken(brCond_io_taken)
  );
  assign io_icache_req_valid = ~stall; // @[Datapath.scala 83:30]
  assign io_icache_req_bits_addr = npc[31:0]; // @[Datapath.scala 80:27]
  assign io_dcache_abort = csr_io__expt | csr_io__vmSwitch; // @[Datapath.scala 200:34]
  assign io_dcache_req_valid = _T_24 & (|io_ctrl_st_type | |io_ctrl_ld_type); // @[Datapath.scala 127:37]
  assign io_dcache_req_bits_addr = daddr[31:0]; // @[Datapath.scala 128:27]
  assign io_dcache_req_bits_data = _T_51[31:0]; // @[Datapath.scala 129:27]
  assign io_dcache_req_bits_mask = _T_62[3:0]; // @[Datapath.scala 130:27]
  assign io_ctrl_inst = fe_inst; // @[Datapath.scala 94:17]
  assign io_table_w_data_valid = io_ctrl_dfc_cmd == 3'h1 & ~csr_io__dfc_full & _T_24; // @[Datapath.scala 203:75]
  assign io_table_w_data_bits_listenAddr = _T_32 & rs2hazard ? ew_alu : regFile_io_rdata2; // @[Datapath.scala 112:16]
  assign io_table_w_data_bits_wPid = rs1[15:0]; // @[Datapath.scala 205:29]
  assign io_table_l_data_valid = io_ctrl_dfc_cmd == 3'h2 & _T_24; // @[Datapath.scala 206:55]
  assign io_table_l_data_bits_listenAddr = _T_32 & rs2hazard ? ew_alu : regFile_io_rdata2; // @[Datapath.scala 112:16]
  assign io_table_e_data_ready = ~stall; // @[Datapath.scala 184:28]
  assign io_vmSwitch = csr_io_vmSwitch;
  assign io_in = csr_io_in;
  assign clearPageFault = csr_clearPageFault_0;
  assign satp = csr_satp_0;
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io__stall = ~io_icache_resp_valid | ~io_dcache_resp_valid; // @[Datapath.scala 63:37]
  assign csr_io__cmd = csr_cmd; // @[Datapath.scala 173:19]
  assign csr_io__in = csr_in; // @[Datapath.scala 172:19]
  assign csr_io__pc = ew_pc[31:0]; // @[Datapath.scala 175:19]
  assign csr_io__addr = ew_alu; // @[Datapath.scala 176:19]
  assign csr_io__inst = ew_inst; // @[Datapath.scala 174:19]
  assign csr_io__illegal = illegal; // @[Datapath.scala 177:19]
  assign csr_io__st_type = st_type; // @[Datapath.scala 180:19]
  assign csr_io__ld_type = ld_type; // @[Datapath.scala 179:19]
  assign csr_io__pc_check = pc_check; // @[Datapath.scala 178:19]
  assign csr_io__dfc_cmd = csr_dfc_cmd; // @[Datapath.scala 183:21]
  assign csr_io__dfc_pid = io_table_e_data_valid ? io_table_e_data_bits_pid : 16'h0; // @[Datapath.scala 185:27]
  assign csr_io__table_f_data_valid = io_table_f_data_valid; // @[Datapath.scala 187:18]
  assign csr_io__table_f_data_bits_full_sig = io_table_f_data_bits_full_sig; // @[Datapath.scala 187:18]
  assign csr_uartRxValid_0 = io_rxChannel_valid;
  assign csr_dmmu = pageFault;
  assign csr_immu = pageFault_0;
  assign regFile_clock = clock;
  assign regFile_io_raddr1 = fe_inst[19:15]; // @[Datapath.scala 98:25]
  assign regFile_io_raddr2 = fe_inst[24:20]; // @[Datapath.scala 99:25]
  assign regFile_io_wen = wb_en & _T_24 & _T_71 & _T_73; // @[Datapath.scala 195:56]
  assign regFile_io_waddr = ew_inst[11:7]; // @[Datapath.scala 108:27]
  assign regFile_io_wdata = regWrite[31:0]; // @[Datapath.scala 197:20]
  assign alu_io_A = _T_37[31:0]; // @[Datapath.scala 115:12]
  assign alu_io_B = io_ctrl_B_sel ? rs2 : immGen_io_out; // @[Datapath.scala 116:18]
  assign alu_io_alu_op = io_ctrl_alu_op; // @[Datapath.scala 117:17]
  assign immGen_io_inst = fe_inst; // @[Datapath.scala 104:18]
  assign immGen_io_sel = io_ctrl_imm_sel; // @[Datapath.scala 105:18]
  assign brCond_io_rs1 = wb_sel == 2'h0 & rs1hazard ? ew_alu : regFile_io_rdata1; // @[Datapath.scala 111:16]
  assign brCond_io_rs2 = _T_32 & rs2hazard ? ew_alu : regFile_io_rdata2; // @[Datapath.scala 112:16]
  assign brCond_io_br_type = io_ctrl_br_type; // @[Datapath.scala 122:21]
  always @(posedge clock) begin
    if (reset) begin // @[Datapath.scala 40:24]
      fe_inst <= 32'h13; // @[Datapath.scala 40:24]
    end else if (_T_24) begin // @[Datapath.scala 87:17]
      if (started | io_ctrl_inst_kill | brCond_io_taken | csr_io__expt | csr_io__vmSwitch) begin // @[Datapath.scala 78:17]
        fe_inst <= 32'h13;
      end else begin
        fe_inst <= io_icache_resp_bits_data;
      end
    end
    if (_T_24) begin // @[Datapath.scala 87:17]
      fe_pc <= pc; // @[Datapath.scala 88:13]
    end
    if (reset) begin // @[Datapath.scala 44:24]
      ew_inst <= 32'h13; // @[Datapath.scala 44:24]
    end else if (!(reset | _T_24 & csr_io__expt | _T_24 & csr_io__vmSwitch)) begin // @[Datapath.scala 138:76]
      if (_T_24 & ~csr_io__expt & ~csr_io__vmSwitch) begin // @[Datapath.scala 147:58]
        ew_inst <= fe_inst; // @[Datapath.scala 149:15]
      end
    end
    if (!(reset | _T_24 & csr_io__expt | _T_24 & csr_io__vmSwitch)) begin // @[Datapath.scala 138:76]
      if (_T_24 & ~csr_io__expt & ~csr_io__vmSwitch) begin // @[Datapath.scala 147:58]
        ew_pc <= fe_pc; // @[Datapath.scala 148:15]
      end
    end
    if (!(reset | _T_24 & csr_io__expt | _T_24 & csr_io__vmSwitch)) begin // @[Datapath.scala 138:76]
      if (_T_24 & ~csr_io__expt & ~csr_io__vmSwitch) begin // @[Datapath.scala 147:58]
        ew_alu <= alu_io_out; // @[Datapath.scala 150:15]
      end
    end
    if (!(reset | _T_24 & csr_io__expt | _T_24 & csr_io__vmSwitch)) begin // @[Datapath.scala 138:76]
      if (_T_24 & ~csr_io__expt & ~csr_io__vmSwitch) begin // @[Datapath.scala 147:58]
        if (io_ctrl_imm_sel == 3'h6) begin // @[Datapath.scala 151:21]
          csr_in <= immGen_io_out;
        end else if (wb_sel == 2'h0 & rs1hazard) begin // @[Datapath.scala 111:16]
          csr_in <= ew_alu;
        end else begin
          csr_in <= regFile_io_rdata1;
        end
      end
    end
    if (reset | _T_24 & csr_io__expt | _T_24 & csr_io__vmSwitch) begin // @[Datapath.scala 138:76]
      st_type <= 2'h0; // @[Datapath.scala 139:15]
    end else if (_T_24 & ~csr_io__expt & ~csr_io__vmSwitch) begin // @[Datapath.scala 147:58]
      st_type <= io_ctrl_st_type; // @[Datapath.scala 152:15]
    end
    if (reset | _T_24 & csr_io__expt | _T_24 & csr_io__vmSwitch) begin // @[Datapath.scala 138:76]
      ld_type <= 3'h0; // @[Datapath.scala 140:15]
    end else if (_T_24 & ~csr_io__expt & ~csr_io__vmSwitch) begin // @[Datapath.scala 147:58]
      ld_type <= io_ctrl_ld_type; // @[Datapath.scala 153:15]
    end
    if (!(reset | _T_24 & csr_io__expt | _T_24 & csr_io__vmSwitch)) begin // @[Datapath.scala 138:76]
      if (_T_24 & ~csr_io__expt & ~csr_io__vmSwitch) begin // @[Datapath.scala 147:58]
        wb_sel <= io_ctrl_wb_sel; // @[Datapath.scala 154:15]
      end
    end
    if (reset | _T_24 & csr_io__expt | _T_24 & csr_io__vmSwitch) begin // @[Datapath.scala 138:76]
      wb_en <= 1'h0; // @[Datapath.scala 141:15]
    end else if (_T_24 & ~csr_io__expt & ~csr_io__vmSwitch) begin // @[Datapath.scala 147:58]
      wb_en <= io_ctrl_wb_en; // @[Datapath.scala 155:15]
    end
    if (reset | _T_24 & csr_io__expt | _T_24 & csr_io__vmSwitch) begin // @[Datapath.scala 138:76]
      csr_cmd <= 3'h0; // @[Datapath.scala 142:15]
    end else if (_T_24 & ~csr_io__expt & ~csr_io__vmSwitch) begin // @[Datapath.scala 147:58]
      csr_cmd <= io_ctrl_csr_cmd; // @[Datapath.scala 156:15]
    end
    if (reset | _T_24 & csr_io__expt | _T_24 & csr_io__vmSwitch) begin // @[Datapath.scala 138:76]
      illegal <= 1'h0; // @[Datapath.scala 143:15]
    end else if (_T_24 & ~csr_io__expt & ~csr_io__vmSwitch) begin // @[Datapath.scala 147:58]
      illegal <= io_ctrl_illegal; // @[Datapath.scala 157:15]
    end
    if (reset | _T_24 & csr_io__expt | _T_24 & csr_io__vmSwitch) begin // @[Datapath.scala 138:76]
      pc_check <= 1'h0; // @[Datapath.scala 144:15]
    end else if (_T_24 & ~csr_io__expt & ~csr_io__vmSwitch) begin // @[Datapath.scala 147:58]
      pc_check <= _T_6; // @[Datapath.scala 158:15]
    end
    if (reset | _T_24 & csr_io__expt | _T_24 & csr_io__vmSwitch) begin // @[Datapath.scala 138:76]
      csr_dfc_cmd <= 3'h0; // @[Datapath.scala 146:17]
    end else if (_T_24 & ~csr_io__expt & ~csr_io__vmSwitch) begin // @[Datapath.scala 147:58]
      csr_dfc_cmd <= io_ctrl_dfc_cmd; // @[Datapath.scala 160:17]
    end
    started <= reset; // @[Datapath.scala 62:31]
    if (reset) begin // @[Datapath.scala 64:21]
      pc <= {{1'd0}, _T_4}; // @[Datapath.scala 64:21]
    end else if (!(stall)) begin // @[Datapath.scala 66:17]
      if (csr_io__expt) begin // @[Datapath.scala 66:32]
        pc <= {{1'd0}, csr_io__evec};
      end else if (io_ctrl_pc_sel == 2'h3) begin // @[Datapath.scala 68:17]
        pc <= {{1'd0}, csr_io__epc};
      end else begin
        pc <= _T_17;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fe_inst = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  fe_pc = _RAND_1[32:0];
  _RAND_2 = {1{`RANDOM}};
  ew_inst = _RAND_2[31:0];
  _RAND_3 = {2{`RANDOM}};
  ew_pc = _RAND_3[32:0];
  _RAND_4 = {1{`RANDOM}};
  ew_alu = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  csr_in = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  st_type = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  ld_type = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  wb_sel = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  wb_en = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  csr_cmd = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  illegal = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  pc_check = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  csr_dfc_cmd = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  started = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  pc = _RAND_15[32:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Control(
  input  [31:0] io_inst,
  output [1:0]  io_pc_sel,
  output        io_inst_kill,
  output        io_A_sel,
  output        io_B_sel,
  output [2:0]  io_imm_sel,
  output [3:0]  io_alu_op,
  output [2:0]  io_br_type,
  output [1:0]  io_st_type,
  output [2:0]  io_ld_type,
  output [1:0]  io_wb_sel,
  output        io_wb_en,
  output [2:0]  io_csr_cmd,
  output        io_illegal,
  output [2:0]  io_dfc_cmd
);
  wire [31:0] _T = io_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _T_1 = 32'h37 == _T; // @[Lookup.scala 31:38]
  wire  _T_3 = 32'h17 == _T; // @[Lookup.scala 31:38]
  wire  _T_5 = 32'h6f == _T; // @[Lookup.scala 31:38]
  wire [31:0] _T_6 = io_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _T_7 = 32'h67 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_9 = 32'h63 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_11 = 32'h1063 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_13 = 32'h4063 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_15 = 32'h5063 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_17 = 32'h6063 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_19 = 32'h7063 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_21 = 32'h3 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_23 = 32'h1003 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_25 = 32'h2003 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_27 = 32'h4003 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_29 = 32'h5003 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_31 = 32'h23 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_33 = 32'h1023 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_35 = 32'h2023 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_37 = 32'h13 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_39 = 32'h2013 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_41 = 32'h3013 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_43 = 32'h4013 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_45 = 32'h6013 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_47 = 32'h7013 == _T_6; // @[Lookup.scala 31:38]
  wire [31:0] _T_48 = io_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _T_49 = 32'h1013 == _T_48; // @[Lookup.scala 31:38]
  wire  _T_51 = 32'h5013 == _T_48; // @[Lookup.scala 31:38]
  wire  _T_53 = 32'h40005013 == _T_48; // @[Lookup.scala 31:38]
  wire  _T_55 = 32'h33 == _T_48; // @[Lookup.scala 31:38]
  wire  _T_57 = 32'h40000033 == _T_48; // @[Lookup.scala 31:38]
  wire  _T_59 = 32'h1033 == _T_48; // @[Lookup.scala 31:38]
  wire  _T_61 = 32'h2033 == _T_48; // @[Lookup.scala 31:38]
  wire  _T_63 = 32'h3033 == _T_48; // @[Lookup.scala 31:38]
  wire  _T_65 = 32'h4033 == _T_48; // @[Lookup.scala 31:38]
  wire  _T_67 = 32'h5033 == _T_48; // @[Lookup.scala 31:38]
  wire  _T_69 = 32'h40005033 == _T_48; // @[Lookup.scala 31:38]
  wire  _T_71 = 32'h6033 == _T_48; // @[Lookup.scala 31:38]
  wire  _T_73 = 32'h7033 == _T_48; // @[Lookup.scala 31:38]
  wire [31:0] _T_74 = io_inst & 32'hf00fffff; // @[Lookup.scala 31:38]
  wire  _T_75 = 32'hf == _T_74; // @[Lookup.scala 31:38]
  wire  _T_77 = 32'h100f == io_inst; // @[Lookup.scala 31:38]
  wire  _T_79 = 32'h1073 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_81 = 32'h2073 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_83 = 32'h3073 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_85 = 32'h5073 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_87 = 32'h6073 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_89 = 32'h7073 == _T_6; // @[Lookup.scala 31:38]
  wire  _T_91 = 32'h73 == io_inst; // @[Lookup.scala 31:38]
  wire  _T_93 = 32'h100073 == io_inst; // @[Lookup.scala 31:38]
  wire  _T_95 = 32'h10000073 == io_inst; // @[Lookup.scala 31:38]
  wire  _T_97 = 32'h10200073 == io_inst; // @[Lookup.scala 31:38]
  wire [31:0] _T_98 = io_inst & 32'hfe007fff; // @[Lookup.scala 31:38]
  wire  _T_99 = 32'h74 == _T_98; // @[Lookup.scala 31:38]
  wire [31:0] _T_100 = io_inst & 32'hfe0fffff; // @[Lookup.scala 31:38]
  wire  _T_101 = 32'h75 == _T_100; // @[Lookup.scala 31:38]
  wire [1:0] _T_105 = _T_95 ? 2'h3 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _T_106 = _T_93 ? 2'h0 : _T_105; // @[Lookup.scala 33:37]
  wire [1:0] _T_107 = _T_91 ? 2'h0 : _T_106; // @[Lookup.scala 33:37]
  wire [1:0] _T_108 = _T_89 ? 2'h2 : _T_107; // @[Lookup.scala 33:37]
  wire [1:0] _T_109 = _T_87 ? 2'h2 : _T_108; // @[Lookup.scala 33:37]
  wire [1:0] _T_110 = _T_85 ? 2'h2 : _T_109; // @[Lookup.scala 33:37]
  wire [1:0] _T_111 = _T_83 ? 2'h2 : _T_110; // @[Lookup.scala 33:37]
  wire [1:0] _T_112 = _T_81 ? 2'h2 : _T_111; // @[Lookup.scala 33:37]
  wire [1:0] _T_113 = _T_79 ? 2'h2 : _T_112; // @[Lookup.scala 33:37]
  wire [1:0] _T_114 = _T_77 ? 2'h2 : _T_113; // @[Lookup.scala 33:37]
  wire [1:0] _T_115 = _T_75 ? 2'h0 : _T_114; // @[Lookup.scala 33:37]
  wire [1:0] _T_116 = _T_73 ? 2'h0 : _T_115; // @[Lookup.scala 33:37]
  wire [1:0] _T_117 = _T_71 ? 2'h0 : _T_116; // @[Lookup.scala 33:37]
  wire [1:0] _T_118 = _T_69 ? 2'h0 : _T_117; // @[Lookup.scala 33:37]
  wire [1:0] _T_119 = _T_67 ? 2'h0 : _T_118; // @[Lookup.scala 33:37]
  wire [1:0] _T_120 = _T_65 ? 2'h0 : _T_119; // @[Lookup.scala 33:37]
  wire [1:0] _T_121 = _T_63 ? 2'h0 : _T_120; // @[Lookup.scala 33:37]
  wire [1:0] _T_122 = _T_61 ? 2'h0 : _T_121; // @[Lookup.scala 33:37]
  wire [1:0] _T_123 = _T_59 ? 2'h0 : _T_122; // @[Lookup.scala 33:37]
  wire [1:0] _T_124 = _T_57 ? 2'h0 : _T_123; // @[Lookup.scala 33:37]
  wire [1:0] _T_125 = _T_55 ? 2'h0 : _T_124; // @[Lookup.scala 33:37]
  wire [1:0] _T_126 = _T_53 ? 2'h0 : _T_125; // @[Lookup.scala 33:37]
  wire [1:0] _T_127 = _T_51 ? 2'h0 : _T_126; // @[Lookup.scala 33:37]
  wire [1:0] _T_128 = _T_49 ? 2'h0 : _T_127; // @[Lookup.scala 33:37]
  wire [1:0] _T_129 = _T_47 ? 2'h0 : _T_128; // @[Lookup.scala 33:37]
  wire [1:0] _T_130 = _T_45 ? 2'h0 : _T_129; // @[Lookup.scala 33:37]
  wire [1:0] _T_131 = _T_43 ? 2'h0 : _T_130; // @[Lookup.scala 33:37]
  wire [1:0] _T_132 = _T_41 ? 2'h0 : _T_131; // @[Lookup.scala 33:37]
  wire [1:0] _T_133 = _T_39 ? 2'h0 : _T_132; // @[Lookup.scala 33:37]
  wire [1:0] _T_134 = _T_37 ? 2'h0 : _T_133; // @[Lookup.scala 33:37]
  wire [1:0] _T_135 = _T_35 ? 2'h0 : _T_134; // @[Lookup.scala 33:37]
  wire [1:0] _T_136 = _T_33 ? 2'h0 : _T_135; // @[Lookup.scala 33:37]
  wire [1:0] _T_137 = _T_31 ? 2'h0 : _T_136; // @[Lookup.scala 33:37]
  wire [1:0] _T_138 = _T_29 ? 2'h2 : _T_137; // @[Lookup.scala 33:37]
  wire [1:0] _T_139 = _T_27 ? 2'h2 : _T_138; // @[Lookup.scala 33:37]
  wire [1:0] _T_140 = _T_25 ? 2'h2 : _T_139; // @[Lookup.scala 33:37]
  wire [1:0] _T_141 = _T_23 ? 2'h2 : _T_140; // @[Lookup.scala 33:37]
  wire [1:0] _T_142 = _T_21 ? 2'h2 : _T_141; // @[Lookup.scala 33:37]
  wire [1:0] _T_143 = _T_19 ? 2'h0 : _T_142; // @[Lookup.scala 33:37]
  wire [1:0] _T_144 = _T_17 ? 2'h0 : _T_143; // @[Lookup.scala 33:37]
  wire [1:0] _T_145 = _T_15 ? 2'h0 : _T_144; // @[Lookup.scala 33:37]
  wire [1:0] _T_146 = _T_13 ? 2'h0 : _T_145; // @[Lookup.scala 33:37]
  wire [1:0] _T_147 = _T_11 ? 2'h0 : _T_146; // @[Lookup.scala 33:37]
  wire [1:0] _T_148 = _T_9 ? 2'h0 : _T_147; // @[Lookup.scala 33:37]
  wire [1:0] _T_149 = _T_7 ? 2'h1 : _T_148; // @[Lookup.scala 33:37]
  wire [1:0] _T_150 = _T_5 ? 2'h1 : _T_149; // @[Lookup.scala 33:37]
  wire [1:0] _T_151 = _T_3 ? 2'h0 : _T_150; // @[Lookup.scala 33:37]
  wire  _T_154 = _T_97 ? 1'h0 : _T_99 | _T_101; // @[Lookup.scala 33:37]
  wire  _T_155 = _T_95 ? 1'h0 : _T_154; // @[Lookup.scala 33:37]
  wire  _T_156 = _T_93 ? 1'h0 : _T_155; // @[Lookup.scala 33:37]
  wire  _T_157 = _T_91 ? 1'h0 : _T_156; // @[Lookup.scala 33:37]
  wire  _T_158 = _T_89 ? 1'h0 : _T_157; // @[Lookup.scala 33:37]
  wire  _T_159 = _T_87 ? 1'h0 : _T_158; // @[Lookup.scala 33:37]
  wire  _T_160 = _T_85 ? 1'h0 : _T_159; // @[Lookup.scala 33:37]
  wire  _T_164 = _T_77 ? 1'h0 : _T_79 | (_T_81 | (_T_83 | _T_160)); // @[Lookup.scala 33:37]
  wire  _T_165 = _T_75 ? 1'h0 : _T_164; // @[Lookup.scala 33:37]
  wire  _T_193 = _T_19 ? 1'h0 : _T_21 | (_T_23 | (_T_25 | (_T_27 | (_T_29 | (_T_31 | (_T_33 | (_T_35 | (_T_37 | (_T_39
     | (_T_41 | (_T_43 | (_T_45 | (_T_47 | (_T_49 | (_T_51 | (_T_53 | (_T_55 | (_T_57 | (_T_59 | (_T_61 | (_T_63 | (
    _T_65 | (_T_67 | (_T_69 | (_T_71 | (_T_73 | _T_165)))))))))))))))))))))))))); // @[Lookup.scala 33:37]
  wire  _T_194 = _T_17 ? 1'h0 : _T_193; // @[Lookup.scala 33:37]
  wire  _T_195 = _T_15 ? 1'h0 : _T_194; // @[Lookup.scala 33:37]
  wire  _T_196 = _T_13 ? 1'h0 : _T_195; // @[Lookup.scala 33:37]
  wire  _T_197 = _T_11 ? 1'h0 : _T_196; // @[Lookup.scala 33:37]
  wire  _T_198 = _T_9 ? 1'h0 : _T_197; // @[Lookup.scala 33:37]
  wire  _T_200 = _T_5 ? 1'h0 : _T_7 | _T_198; // @[Lookup.scala 33:37]
  wire  _T_201 = _T_3 ? 1'h0 : _T_200; // @[Lookup.scala 33:37]
  wire  _T_204 = _T_97 ? 1'h0 : _T_99; // @[Lookup.scala 33:37]
  wire  _T_205 = _T_95 ? 1'h0 : _T_204; // @[Lookup.scala 33:37]
  wire  _T_206 = _T_93 ? 1'h0 : _T_205; // @[Lookup.scala 33:37]
  wire  _T_207 = _T_91 ? 1'h0 : _T_206; // @[Lookup.scala 33:37]
  wire  _T_208 = _T_89 ? 1'h0 : _T_207; // @[Lookup.scala 33:37]
  wire  _T_209 = _T_87 ? 1'h0 : _T_208; // @[Lookup.scala 33:37]
  wire  _T_210 = _T_85 ? 1'h0 : _T_209; // @[Lookup.scala 33:37]
  wire  _T_211 = _T_83 ? 1'h0 : _T_210; // @[Lookup.scala 33:37]
  wire  _T_212 = _T_81 ? 1'h0 : _T_211; // @[Lookup.scala 33:37]
  wire  _T_213 = _T_79 ? 1'h0 : _T_212; // @[Lookup.scala 33:37]
  wire  _T_214 = _T_77 ? 1'h0 : _T_213; // @[Lookup.scala 33:37]
  wire  _T_215 = _T_75 ? 1'h0 : _T_214; // @[Lookup.scala 33:37]
  wire  _T_226 = _T_53 ? 1'h0 : _T_55 | (_T_57 | (_T_59 | (_T_61 | (_T_63 | (_T_65 | (_T_67 | (_T_69 | (_T_71 | (_T_73
     | _T_215))))))))); // @[Lookup.scala 33:37]
  wire  _T_227 = _T_51 ? 1'h0 : _T_226; // @[Lookup.scala 33:37]
  wire  _T_228 = _T_49 ? 1'h0 : _T_227; // @[Lookup.scala 33:37]
  wire  _T_229 = _T_47 ? 1'h0 : _T_228; // @[Lookup.scala 33:37]
  wire  _T_230 = _T_45 ? 1'h0 : _T_229; // @[Lookup.scala 33:37]
  wire  _T_231 = _T_43 ? 1'h0 : _T_230; // @[Lookup.scala 33:37]
  wire  _T_232 = _T_41 ? 1'h0 : _T_231; // @[Lookup.scala 33:37]
  wire  _T_233 = _T_39 ? 1'h0 : _T_232; // @[Lookup.scala 33:37]
  wire  _T_234 = _T_37 ? 1'h0 : _T_233; // @[Lookup.scala 33:37]
  wire  _T_235 = _T_35 ? 1'h0 : _T_234; // @[Lookup.scala 33:37]
  wire  _T_236 = _T_33 ? 1'h0 : _T_235; // @[Lookup.scala 33:37]
  wire  _T_237 = _T_31 ? 1'h0 : _T_236; // @[Lookup.scala 33:37]
  wire  _T_238 = _T_29 ? 1'h0 : _T_237; // @[Lookup.scala 33:37]
  wire  _T_239 = _T_27 ? 1'h0 : _T_238; // @[Lookup.scala 33:37]
  wire  _T_240 = _T_25 ? 1'h0 : _T_239; // @[Lookup.scala 33:37]
  wire  _T_241 = _T_23 ? 1'h0 : _T_240; // @[Lookup.scala 33:37]
  wire  _T_242 = _T_21 ? 1'h0 : _T_241; // @[Lookup.scala 33:37]
  wire  _T_243 = _T_19 ? 1'h0 : _T_242; // @[Lookup.scala 33:37]
  wire  _T_244 = _T_17 ? 1'h0 : _T_243; // @[Lookup.scala 33:37]
  wire  _T_245 = _T_15 ? 1'h0 : _T_244; // @[Lookup.scala 33:37]
  wire  _T_246 = _T_13 ? 1'h0 : _T_245; // @[Lookup.scala 33:37]
  wire  _T_247 = _T_11 ? 1'h0 : _T_246; // @[Lookup.scala 33:37]
  wire  _T_248 = _T_9 ? 1'h0 : _T_247; // @[Lookup.scala 33:37]
  wire  _T_249 = _T_7 ? 1'h0 : _T_248; // @[Lookup.scala 33:37]
  wire  _T_250 = _T_5 ? 1'h0 : _T_249; // @[Lookup.scala 33:37]
  wire  _T_251 = _T_3 ? 1'h0 : _T_250; // @[Lookup.scala 33:37]
  wire [2:0] _T_258 = _T_89 ? 3'h6 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_259 = _T_87 ? 3'h6 : _T_258; // @[Lookup.scala 33:37]
  wire [2:0] _T_260 = _T_85 ? 3'h6 : _T_259; // @[Lookup.scala 33:37]
  wire [2:0] _T_261 = _T_83 ? 3'h0 : _T_260; // @[Lookup.scala 33:37]
  wire [2:0] _T_262 = _T_81 ? 3'h0 : _T_261; // @[Lookup.scala 33:37]
  wire [2:0] _T_263 = _T_79 ? 3'h0 : _T_262; // @[Lookup.scala 33:37]
  wire [2:0] _T_264 = _T_77 ? 3'h0 : _T_263; // @[Lookup.scala 33:37]
  wire [2:0] _T_265 = _T_75 ? 3'h0 : _T_264; // @[Lookup.scala 33:37]
  wire [2:0] _T_266 = _T_73 ? 3'h0 : _T_265; // @[Lookup.scala 33:37]
  wire [2:0] _T_267 = _T_71 ? 3'h0 : _T_266; // @[Lookup.scala 33:37]
  wire [2:0] _T_268 = _T_69 ? 3'h0 : _T_267; // @[Lookup.scala 33:37]
  wire [2:0] _T_269 = _T_67 ? 3'h0 : _T_268; // @[Lookup.scala 33:37]
  wire [2:0] _T_270 = _T_65 ? 3'h0 : _T_269; // @[Lookup.scala 33:37]
  wire [2:0] _T_271 = _T_63 ? 3'h0 : _T_270; // @[Lookup.scala 33:37]
  wire [2:0] _T_272 = _T_61 ? 3'h0 : _T_271; // @[Lookup.scala 33:37]
  wire [2:0] _T_273 = _T_59 ? 3'h0 : _T_272; // @[Lookup.scala 33:37]
  wire [2:0] _T_274 = _T_57 ? 3'h0 : _T_273; // @[Lookup.scala 33:37]
  wire [2:0] _T_275 = _T_55 ? 3'h0 : _T_274; // @[Lookup.scala 33:37]
  wire [2:0] _T_276 = _T_53 ? 3'h1 : _T_275; // @[Lookup.scala 33:37]
  wire [2:0] _T_277 = _T_51 ? 3'h1 : _T_276; // @[Lookup.scala 33:37]
  wire [2:0] _T_278 = _T_49 ? 3'h1 : _T_277; // @[Lookup.scala 33:37]
  wire [2:0] _T_279 = _T_47 ? 3'h1 : _T_278; // @[Lookup.scala 33:37]
  wire [2:0] _T_280 = _T_45 ? 3'h1 : _T_279; // @[Lookup.scala 33:37]
  wire [2:0] _T_281 = _T_43 ? 3'h1 : _T_280; // @[Lookup.scala 33:37]
  wire [2:0] _T_282 = _T_41 ? 3'h1 : _T_281; // @[Lookup.scala 33:37]
  wire [2:0] _T_283 = _T_39 ? 3'h1 : _T_282; // @[Lookup.scala 33:37]
  wire [2:0] _T_284 = _T_37 ? 3'h1 : _T_283; // @[Lookup.scala 33:37]
  wire [2:0] _T_285 = _T_35 ? 3'h2 : _T_284; // @[Lookup.scala 33:37]
  wire [2:0] _T_286 = _T_33 ? 3'h2 : _T_285; // @[Lookup.scala 33:37]
  wire [2:0] _T_287 = _T_31 ? 3'h2 : _T_286; // @[Lookup.scala 33:37]
  wire [2:0] _T_288 = _T_29 ? 3'h1 : _T_287; // @[Lookup.scala 33:37]
  wire [2:0] _T_289 = _T_27 ? 3'h1 : _T_288; // @[Lookup.scala 33:37]
  wire [2:0] _T_290 = _T_25 ? 3'h1 : _T_289; // @[Lookup.scala 33:37]
  wire [2:0] _T_291 = _T_23 ? 3'h1 : _T_290; // @[Lookup.scala 33:37]
  wire [2:0] _T_292 = _T_21 ? 3'h1 : _T_291; // @[Lookup.scala 33:37]
  wire [2:0] _T_293 = _T_19 ? 3'h5 : _T_292; // @[Lookup.scala 33:37]
  wire [2:0] _T_294 = _T_17 ? 3'h5 : _T_293; // @[Lookup.scala 33:37]
  wire [2:0] _T_295 = _T_15 ? 3'h5 : _T_294; // @[Lookup.scala 33:37]
  wire [2:0] _T_296 = _T_13 ? 3'h5 : _T_295; // @[Lookup.scala 33:37]
  wire [2:0] _T_297 = _T_11 ? 3'h5 : _T_296; // @[Lookup.scala 33:37]
  wire [2:0] _T_298 = _T_9 ? 3'h5 : _T_297; // @[Lookup.scala 33:37]
  wire [2:0] _T_299 = _T_7 ? 3'h1 : _T_298; // @[Lookup.scala 33:37]
  wire [2:0] _T_300 = _T_5 ? 3'h4 : _T_299; // @[Lookup.scala 33:37]
  wire [2:0] _T_301 = _T_3 ? 3'h3 : _T_300; // @[Lookup.scala 33:37]
  wire [3:0] _T_311 = _T_83 ? 4'ha : 4'hf; // @[Lookup.scala 33:37]
  wire [3:0] _T_312 = _T_81 ? 4'ha : _T_311; // @[Lookup.scala 33:37]
  wire [3:0] _T_313 = _T_79 ? 4'ha : _T_312; // @[Lookup.scala 33:37]
  wire [3:0] _T_314 = _T_77 ? 4'hf : _T_313; // @[Lookup.scala 33:37]
  wire [3:0] _T_315 = _T_75 ? 4'hf : _T_314; // @[Lookup.scala 33:37]
  wire [3:0] _T_316 = _T_73 ? 4'h2 : _T_315; // @[Lookup.scala 33:37]
  wire [3:0] _T_317 = _T_71 ? 4'h3 : _T_316; // @[Lookup.scala 33:37]
  wire [3:0] _T_318 = _T_69 ? 4'h9 : _T_317; // @[Lookup.scala 33:37]
  wire [3:0] _T_319 = _T_67 ? 4'h8 : _T_318; // @[Lookup.scala 33:37]
  wire [3:0] _T_320 = _T_65 ? 4'h4 : _T_319; // @[Lookup.scala 33:37]
  wire [3:0] _T_321 = _T_63 ? 4'h7 : _T_320; // @[Lookup.scala 33:37]
  wire [3:0] _T_322 = _T_61 ? 4'h5 : _T_321; // @[Lookup.scala 33:37]
  wire [3:0] _T_323 = _T_59 ? 4'h6 : _T_322; // @[Lookup.scala 33:37]
  wire [3:0] _T_324 = _T_57 ? 4'h1 : _T_323; // @[Lookup.scala 33:37]
  wire [3:0] _T_325 = _T_55 ? 4'h0 : _T_324; // @[Lookup.scala 33:37]
  wire [3:0] _T_326 = _T_53 ? 4'h9 : _T_325; // @[Lookup.scala 33:37]
  wire [3:0] _T_327 = _T_51 ? 4'h8 : _T_326; // @[Lookup.scala 33:37]
  wire [3:0] _T_328 = _T_49 ? 4'h6 : _T_327; // @[Lookup.scala 33:37]
  wire [3:0] _T_329 = _T_47 ? 4'h2 : _T_328; // @[Lookup.scala 33:37]
  wire [3:0] _T_330 = _T_45 ? 4'h3 : _T_329; // @[Lookup.scala 33:37]
  wire [3:0] _T_331 = _T_43 ? 4'h4 : _T_330; // @[Lookup.scala 33:37]
  wire [3:0] _T_332 = _T_41 ? 4'h7 : _T_331; // @[Lookup.scala 33:37]
  wire [3:0] _T_333 = _T_39 ? 4'h5 : _T_332; // @[Lookup.scala 33:37]
  wire [3:0] _T_334 = _T_37 ? 4'h0 : _T_333; // @[Lookup.scala 33:37]
  wire [3:0] _T_335 = _T_35 ? 4'h0 : _T_334; // @[Lookup.scala 33:37]
  wire [3:0] _T_336 = _T_33 ? 4'h0 : _T_335; // @[Lookup.scala 33:37]
  wire [3:0] _T_337 = _T_31 ? 4'h0 : _T_336; // @[Lookup.scala 33:37]
  wire [3:0] _T_338 = _T_29 ? 4'h0 : _T_337; // @[Lookup.scala 33:37]
  wire [3:0] _T_339 = _T_27 ? 4'h0 : _T_338; // @[Lookup.scala 33:37]
  wire [3:0] _T_340 = _T_25 ? 4'h0 : _T_339; // @[Lookup.scala 33:37]
  wire [3:0] _T_341 = _T_23 ? 4'h0 : _T_340; // @[Lookup.scala 33:37]
  wire [3:0] _T_342 = _T_21 ? 4'h0 : _T_341; // @[Lookup.scala 33:37]
  wire [3:0] _T_343 = _T_19 ? 4'h0 : _T_342; // @[Lookup.scala 33:37]
  wire [3:0] _T_344 = _T_17 ? 4'h0 : _T_343; // @[Lookup.scala 33:37]
  wire [3:0] _T_345 = _T_15 ? 4'h0 : _T_344; // @[Lookup.scala 33:37]
  wire [3:0] _T_346 = _T_13 ? 4'h0 : _T_345; // @[Lookup.scala 33:37]
  wire [3:0] _T_347 = _T_11 ? 4'h0 : _T_346; // @[Lookup.scala 33:37]
  wire [3:0] _T_348 = _T_9 ? 4'h0 : _T_347; // @[Lookup.scala 33:37]
  wire [3:0] _T_349 = _T_7 ? 4'h0 : _T_348; // @[Lookup.scala 33:37]
  wire [3:0] _T_350 = _T_5 ? 4'h0 : _T_349; // @[Lookup.scala 33:37]
  wire [3:0] _T_351 = _T_3 ? 4'h0 : _T_350; // @[Lookup.scala 33:37]
  wire [2:0] _T_393 = _T_19 ? 3'h4 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_394 = _T_17 ? 3'h1 : _T_393; // @[Lookup.scala 33:37]
  wire [2:0] _T_395 = _T_15 ? 3'h5 : _T_394; // @[Lookup.scala 33:37]
  wire [2:0] _T_396 = _T_13 ? 3'h2 : _T_395; // @[Lookup.scala 33:37]
  wire [2:0] _T_397 = _T_11 ? 3'h6 : _T_396; // @[Lookup.scala 33:37]
  wire [2:0] _T_398 = _T_9 ? 3'h3 : _T_397; // @[Lookup.scala 33:37]
  wire [2:0] _T_399 = _T_7 ? 3'h0 : _T_398; // @[Lookup.scala 33:37]
  wire [2:0] _T_400 = _T_5 ? 3'h0 : _T_399; // @[Lookup.scala 33:37]
  wire [2:0] _T_401 = _T_3 ? 3'h0 : _T_400; // @[Lookup.scala 33:37]
  wire  _T_406 = _T_93 ? 1'h0 : _T_95; // @[Lookup.scala 33:37]
  wire  _T_407 = _T_91 ? 1'h0 : _T_406; // @[Lookup.scala 33:37]
  wire  _T_415 = _T_75 ? 1'h0 : _T_77 | (_T_79 | (_T_81 | (_T_83 | (_T_85 | (_T_87 | (_T_89 | _T_407)))))); // @[Lookup.scala 33:37]
  wire  _T_416 = _T_73 ? 1'h0 : _T_415; // @[Lookup.scala 33:37]
  wire  _T_417 = _T_71 ? 1'h0 : _T_416; // @[Lookup.scala 33:37]
  wire  _T_418 = _T_69 ? 1'h0 : _T_417; // @[Lookup.scala 33:37]
  wire  _T_419 = _T_67 ? 1'h0 : _T_418; // @[Lookup.scala 33:37]
  wire  _T_420 = _T_65 ? 1'h0 : _T_419; // @[Lookup.scala 33:37]
  wire  _T_421 = _T_63 ? 1'h0 : _T_420; // @[Lookup.scala 33:37]
  wire  _T_422 = _T_61 ? 1'h0 : _T_421; // @[Lookup.scala 33:37]
  wire  _T_423 = _T_59 ? 1'h0 : _T_422; // @[Lookup.scala 33:37]
  wire  _T_424 = _T_57 ? 1'h0 : _T_423; // @[Lookup.scala 33:37]
  wire  _T_425 = _T_55 ? 1'h0 : _T_424; // @[Lookup.scala 33:37]
  wire  _T_426 = _T_53 ? 1'h0 : _T_425; // @[Lookup.scala 33:37]
  wire  _T_427 = _T_51 ? 1'h0 : _T_426; // @[Lookup.scala 33:37]
  wire  _T_428 = _T_49 ? 1'h0 : _T_427; // @[Lookup.scala 33:37]
  wire  _T_429 = _T_47 ? 1'h0 : _T_428; // @[Lookup.scala 33:37]
  wire  _T_430 = _T_45 ? 1'h0 : _T_429; // @[Lookup.scala 33:37]
  wire  _T_431 = _T_43 ? 1'h0 : _T_430; // @[Lookup.scala 33:37]
  wire  _T_432 = _T_41 ? 1'h0 : _T_431; // @[Lookup.scala 33:37]
  wire  _T_433 = _T_39 ? 1'h0 : _T_432; // @[Lookup.scala 33:37]
  wire  _T_434 = _T_37 ? 1'h0 : _T_433; // @[Lookup.scala 33:37]
  wire  _T_435 = _T_35 ? 1'h0 : _T_434; // @[Lookup.scala 33:37]
  wire  _T_436 = _T_33 ? 1'h0 : _T_435; // @[Lookup.scala 33:37]
  wire  _T_437 = _T_31 ? 1'h0 : _T_436; // @[Lookup.scala 33:37]
  wire  _T_443 = _T_19 ? 1'h0 : _T_21 | (_T_23 | (_T_25 | (_T_27 | (_T_29 | _T_437)))); // @[Lookup.scala 33:37]
  wire  _T_444 = _T_17 ? 1'h0 : _T_443; // @[Lookup.scala 33:37]
  wire  _T_445 = _T_15 ? 1'h0 : _T_444; // @[Lookup.scala 33:37]
  wire  _T_446 = _T_13 ? 1'h0 : _T_445; // @[Lookup.scala 33:37]
  wire  _T_447 = _T_11 ? 1'h0 : _T_446; // @[Lookup.scala 33:37]
  wire  _T_448 = _T_9 ? 1'h0 : _T_447; // @[Lookup.scala 33:37]
  wire  _T_451 = _T_3 ? 1'h0 : _T_5 | (_T_7 | _T_448); // @[Lookup.scala 33:37]
  wire [1:0] _T_485 = _T_35 ? 2'h1 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _T_486 = _T_33 ? 2'h2 : _T_485; // @[Lookup.scala 33:37]
  wire [1:0] _T_487 = _T_31 ? 2'h3 : _T_486; // @[Lookup.scala 33:37]
  wire [1:0] _T_488 = _T_29 ? 2'h0 : _T_487; // @[Lookup.scala 33:37]
  wire [1:0] _T_489 = _T_27 ? 2'h0 : _T_488; // @[Lookup.scala 33:37]
  wire [1:0] _T_490 = _T_25 ? 2'h0 : _T_489; // @[Lookup.scala 33:37]
  wire [1:0] _T_491 = _T_23 ? 2'h0 : _T_490; // @[Lookup.scala 33:37]
  wire [1:0] _T_492 = _T_21 ? 2'h0 : _T_491; // @[Lookup.scala 33:37]
  wire [1:0] _T_493 = _T_19 ? 2'h0 : _T_492; // @[Lookup.scala 33:37]
  wire [1:0] _T_494 = _T_17 ? 2'h0 : _T_493; // @[Lookup.scala 33:37]
  wire [1:0] _T_495 = _T_15 ? 2'h0 : _T_494; // @[Lookup.scala 33:37]
  wire [1:0] _T_496 = _T_13 ? 2'h0 : _T_495; // @[Lookup.scala 33:37]
  wire [1:0] _T_497 = _T_11 ? 2'h0 : _T_496; // @[Lookup.scala 33:37]
  wire [1:0] _T_498 = _T_9 ? 2'h0 : _T_497; // @[Lookup.scala 33:37]
  wire [1:0] _T_499 = _T_7 ? 2'h0 : _T_498; // @[Lookup.scala 33:37]
  wire [1:0] _T_500 = _T_5 ? 2'h0 : _T_499; // @[Lookup.scala 33:37]
  wire [1:0] _T_501 = _T_3 ? 2'h0 : _T_500; // @[Lookup.scala 33:37]
  wire [2:0] _T_538 = _T_29 ? 3'h4 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_539 = _T_27 ? 3'h5 : _T_538; // @[Lookup.scala 33:37]
  wire [2:0] _T_540 = _T_25 ? 3'h1 : _T_539; // @[Lookup.scala 33:37]
  wire [2:0] _T_541 = _T_23 ? 3'h2 : _T_540; // @[Lookup.scala 33:37]
  wire [2:0] _T_542 = _T_21 ? 3'h3 : _T_541; // @[Lookup.scala 33:37]
  wire [2:0] _T_543 = _T_19 ? 3'h0 : _T_542; // @[Lookup.scala 33:37]
  wire [2:0] _T_544 = _T_17 ? 3'h0 : _T_543; // @[Lookup.scala 33:37]
  wire [2:0] _T_545 = _T_15 ? 3'h0 : _T_544; // @[Lookup.scala 33:37]
  wire [2:0] _T_546 = _T_13 ? 3'h0 : _T_545; // @[Lookup.scala 33:37]
  wire [2:0] _T_547 = _T_11 ? 3'h0 : _T_546; // @[Lookup.scala 33:37]
  wire [2:0] _T_548 = _T_9 ? 3'h0 : _T_547; // @[Lookup.scala 33:37]
  wire [2:0] _T_549 = _T_7 ? 3'h0 : _T_548; // @[Lookup.scala 33:37]
  wire [2:0] _T_550 = _T_5 ? 3'h0 : _T_549; // @[Lookup.scala 33:37]
  wire [2:0] _T_551 = _T_3 ? 3'h0 : _T_550; // @[Lookup.scala 33:37]
  wire [1:0] _T_556 = _T_93 ? 2'h3 : _T_105; // @[Lookup.scala 33:37]
  wire [1:0] _T_557 = _T_91 ? 2'h3 : _T_556; // @[Lookup.scala 33:37]
  wire [1:0] _T_558 = _T_89 ? 2'h3 : _T_557; // @[Lookup.scala 33:37]
  wire [1:0] _T_559 = _T_87 ? 2'h3 : _T_558; // @[Lookup.scala 33:37]
  wire [1:0] _T_560 = _T_85 ? 2'h3 : _T_559; // @[Lookup.scala 33:37]
  wire [1:0] _T_561 = _T_83 ? 2'h3 : _T_560; // @[Lookup.scala 33:37]
  wire [1:0] _T_562 = _T_81 ? 2'h3 : _T_561; // @[Lookup.scala 33:37]
  wire [1:0] _T_563 = _T_79 ? 2'h3 : _T_562; // @[Lookup.scala 33:37]
  wire [1:0] _T_564 = _T_77 ? 2'h0 : _T_563; // @[Lookup.scala 33:37]
  wire [1:0] _T_565 = _T_75 ? 2'h0 : _T_564; // @[Lookup.scala 33:37]
  wire [1:0] _T_566 = _T_73 ? 2'h0 : _T_565; // @[Lookup.scala 33:37]
  wire [1:0] _T_567 = _T_71 ? 2'h0 : _T_566; // @[Lookup.scala 33:37]
  wire [1:0] _T_568 = _T_69 ? 2'h0 : _T_567; // @[Lookup.scala 33:37]
  wire [1:0] _T_569 = _T_67 ? 2'h0 : _T_568; // @[Lookup.scala 33:37]
  wire [1:0] _T_570 = _T_65 ? 2'h0 : _T_569; // @[Lookup.scala 33:37]
  wire [1:0] _T_571 = _T_63 ? 2'h0 : _T_570; // @[Lookup.scala 33:37]
  wire [1:0] _T_572 = _T_61 ? 2'h0 : _T_571; // @[Lookup.scala 33:37]
  wire [1:0] _T_573 = _T_59 ? 2'h0 : _T_572; // @[Lookup.scala 33:37]
  wire [1:0] _T_574 = _T_57 ? 2'h0 : _T_573; // @[Lookup.scala 33:37]
  wire [1:0] _T_575 = _T_55 ? 2'h0 : _T_574; // @[Lookup.scala 33:37]
  wire [1:0] _T_576 = _T_53 ? 2'h0 : _T_575; // @[Lookup.scala 33:37]
  wire [1:0] _T_577 = _T_51 ? 2'h0 : _T_576; // @[Lookup.scala 33:37]
  wire [1:0] _T_578 = _T_49 ? 2'h0 : _T_577; // @[Lookup.scala 33:37]
  wire [1:0] _T_579 = _T_47 ? 2'h0 : _T_578; // @[Lookup.scala 33:37]
  wire [1:0] _T_580 = _T_45 ? 2'h0 : _T_579; // @[Lookup.scala 33:37]
  wire [1:0] _T_581 = _T_43 ? 2'h0 : _T_580; // @[Lookup.scala 33:37]
  wire [1:0] _T_582 = _T_41 ? 2'h0 : _T_581; // @[Lookup.scala 33:37]
  wire [1:0] _T_583 = _T_39 ? 2'h0 : _T_582; // @[Lookup.scala 33:37]
  wire [1:0] _T_584 = _T_37 ? 2'h0 : _T_583; // @[Lookup.scala 33:37]
  wire [1:0] _T_585 = _T_35 ? 2'h0 : _T_584; // @[Lookup.scala 33:37]
  wire [1:0] _T_586 = _T_33 ? 2'h0 : _T_585; // @[Lookup.scala 33:37]
  wire [1:0] _T_587 = _T_31 ? 2'h0 : _T_586; // @[Lookup.scala 33:37]
  wire [1:0] _T_588 = _T_29 ? 2'h1 : _T_587; // @[Lookup.scala 33:37]
  wire [1:0] _T_589 = _T_27 ? 2'h1 : _T_588; // @[Lookup.scala 33:37]
  wire [1:0] _T_590 = _T_25 ? 2'h1 : _T_589; // @[Lookup.scala 33:37]
  wire [1:0] _T_591 = _T_23 ? 2'h1 : _T_590; // @[Lookup.scala 33:37]
  wire [1:0] _T_592 = _T_21 ? 2'h1 : _T_591; // @[Lookup.scala 33:37]
  wire [1:0] _T_593 = _T_19 ? 2'h0 : _T_592; // @[Lookup.scala 33:37]
  wire [1:0] _T_594 = _T_17 ? 2'h0 : _T_593; // @[Lookup.scala 33:37]
  wire [1:0] _T_595 = _T_15 ? 2'h0 : _T_594; // @[Lookup.scala 33:37]
  wire [1:0] _T_596 = _T_13 ? 2'h0 : _T_595; // @[Lookup.scala 33:37]
  wire [1:0] _T_597 = _T_11 ? 2'h0 : _T_596; // @[Lookup.scala 33:37]
  wire [1:0] _T_598 = _T_9 ? 2'h0 : _T_597; // @[Lookup.scala 33:37]
  wire [1:0] _T_599 = _T_7 ? 2'h2 : _T_598; // @[Lookup.scala 33:37]
  wire [1:0] _T_600 = _T_5 ? 2'h2 : _T_599; // @[Lookup.scala 33:37]
  wire [1:0] _T_601 = _T_3 ? 2'h0 : _T_600; // @[Lookup.scala 33:37]
  wire  _T_614 = _T_77 ? 1'h0 : _T_79 | (_T_81 | (_T_83 | (_T_85 | (_T_87 | _T_89)))); // @[Lookup.scala 33:37]
  wire  _T_615 = _T_75 ? 1'h0 : _T_614; // @[Lookup.scala 33:37]
  wire  _T_635 = _T_35 ? 1'h0 : _T_37 | (_T_39 | (_T_41 | (_T_43 | (_T_45 | (_T_47 | (_T_49 | (_T_51 | (_T_53 | (_T_55
     | (_T_57 | (_T_59 | (_T_61 | (_T_63 | (_T_65 | (_T_67 | (_T_69 | (_T_71 | (_T_73 | _T_615)))))))))))))))))); // @[Lookup.scala 33:37]
  wire  _T_636 = _T_33 ? 1'h0 : _T_635; // @[Lookup.scala 33:37]
  wire  _T_637 = _T_31 ? 1'h0 : _T_636; // @[Lookup.scala 33:37]
  wire  _T_643 = _T_19 ? 1'h0 : _T_21 | (_T_23 | (_T_25 | (_T_27 | (_T_29 | _T_637)))); // @[Lookup.scala 33:37]
  wire  _T_644 = _T_17 ? 1'h0 : _T_643; // @[Lookup.scala 33:37]
  wire  _T_645 = _T_15 ? 1'h0 : _T_644; // @[Lookup.scala 33:37]
  wire  _T_646 = _T_13 ? 1'h0 : _T_645; // @[Lookup.scala 33:37]
  wire  _T_647 = _T_11 ? 1'h0 : _T_646; // @[Lookup.scala 33:37]
  wire  _T_648 = _T_9 ? 1'h0 : _T_647; // @[Lookup.scala 33:37]
  wire [2:0] _T_655 = _T_95 ? 3'h4 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_656 = _T_93 ? 3'h4 : _T_655; // @[Lookup.scala 33:37]
  wire [2:0] _T_657 = _T_91 ? 3'h4 : _T_656; // @[Lookup.scala 33:37]
  wire [2:0] _T_658 = _T_89 ? 3'h3 : _T_657; // @[Lookup.scala 33:37]
  wire [2:0] _T_659 = _T_87 ? 3'h2 : _T_658; // @[Lookup.scala 33:37]
  wire [2:0] _T_660 = _T_85 ? 3'h1 : _T_659; // @[Lookup.scala 33:37]
  wire [2:0] _T_661 = _T_83 ? 3'h3 : _T_660; // @[Lookup.scala 33:37]
  wire [2:0] _T_662 = _T_81 ? 3'h2 : _T_661; // @[Lookup.scala 33:37]
  wire [2:0] _T_663 = _T_79 ? 3'h1 : _T_662; // @[Lookup.scala 33:37]
  wire [2:0] _T_664 = _T_77 ? 3'h0 : _T_663; // @[Lookup.scala 33:37]
  wire [2:0] _T_665 = _T_75 ? 3'h0 : _T_664; // @[Lookup.scala 33:37]
  wire [2:0] _T_666 = _T_73 ? 3'h0 : _T_665; // @[Lookup.scala 33:37]
  wire [2:0] _T_667 = _T_71 ? 3'h0 : _T_666; // @[Lookup.scala 33:37]
  wire [2:0] _T_668 = _T_69 ? 3'h0 : _T_667; // @[Lookup.scala 33:37]
  wire [2:0] _T_669 = _T_67 ? 3'h0 : _T_668; // @[Lookup.scala 33:37]
  wire [2:0] _T_670 = _T_65 ? 3'h0 : _T_669; // @[Lookup.scala 33:37]
  wire [2:0] _T_671 = _T_63 ? 3'h0 : _T_670; // @[Lookup.scala 33:37]
  wire [2:0] _T_672 = _T_61 ? 3'h0 : _T_671; // @[Lookup.scala 33:37]
  wire [2:0] _T_673 = _T_59 ? 3'h0 : _T_672; // @[Lookup.scala 33:37]
  wire [2:0] _T_674 = _T_57 ? 3'h0 : _T_673; // @[Lookup.scala 33:37]
  wire [2:0] _T_675 = _T_55 ? 3'h0 : _T_674; // @[Lookup.scala 33:37]
  wire [2:0] _T_676 = _T_53 ? 3'h0 : _T_675; // @[Lookup.scala 33:37]
  wire [2:0] _T_677 = _T_51 ? 3'h0 : _T_676; // @[Lookup.scala 33:37]
  wire [2:0] _T_678 = _T_49 ? 3'h0 : _T_677; // @[Lookup.scala 33:37]
  wire [2:0] _T_679 = _T_47 ? 3'h0 : _T_678; // @[Lookup.scala 33:37]
  wire [2:0] _T_680 = _T_45 ? 3'h0 : _T_679; // @[Lookup.scala 33:37]
  wire [2:0] _T_681 = _T_43 ? 3'h0 : _T_680; // @[Lookup.scala 33:37]
  wire [2:0] _T_682 = _T_41 ? 3'h0 : _T_681; // @[Lookup.scala 33:37]
  wire [2:0] _T_683 = _T_39 ? 3'h0 : _T_682; // @[Lookup.scala 33:37]
  wire [2:0] _T_684 = _T_37 ? 3'h0 : _T_683; // @[Lookup.scala 33:37]
  wire [2:0] _T_685 = _T_35 ? 3'h0 : _T_684; // @[Lookup.scala 33:37]
  wire [2:0] _T_686 = _T_33 ? 3'h0 : _T_685; // @[Lookup.scala 33:37]
  wire [2:0] _T_687 = _T_31 ? 3'h0 : _T_686; // @[Lookup.scala 33:37]
  wire [2:0] _T_688 = _T_29 ? 3'h0 : _T_687; // @[Lookup.scala 33:37]
  wire [2:0] _T_689 = _T_27 ? 3'h0 : _T_688; // @[Lookup.scala 33:37]
  wire [2:0] _T_690 = _T_25 ? 3'h0 : _T_689; // @[Lookup.scala 33:37]
  wire [2:0] _T_691 = _T_23 ? 3'h0 : _T_690; // @[Lookup.scala 33:37]
  wire [2:0] _T_692 = _T_21 ? 3'h0 : _T_691; // @[Lookup.scala 33:37]
  wire [2:0] _T_693 = _T_19 ? 3'h0 : _T_692; // @[Lookup.scala 33:37]
  wire [2:0] _T_694 = _T_17 ? 3'h0 : _T_693; // @[Lookup.scala 33:37]
  wire [2:0] _T_695 = _T_15 ? 3'h0 : _T_694; // @[Lookup.scala 33:37]
  wire [2:0] _T_696 = _T_13 ? 3'h0 : _T_695; // @[Lookup.scala 33:37]
  wire [2:0] _T_697 = _T_11 ? 3'h0 : _T_696; // @[Lookup.scala 33:37]
  wire [2:0] _T_698 = _T_9 ? 3'h0 : _T_697; // @[Lookup.scala 33:37]
  wire [2:0] _T_699 = _T_7 ? 3'h0 : _T_698; // @[Lookup.scala 33:37]
  wire [2:0] _T_700 = _T_5 ? 3'h0 : _T_699; // @[Lookup.scala 33:37]
  wire [2:0] _T_701 = _T_3 ? 3'h0 : _T_700; // @[Lookup.scala 33:37]
  wire  _T_702 = _T_101 ? 1'h0 : 1'h1; // @[Lookup.scala 33:37]
  wire  _T_703 = _T_99 ? 1'h0 : _T_702; // @[Lookup.scala 33:37]
  wire  _T_704 = _T_97 ? 1'h0 : _T_703; // @[Lookup.scala 33:37]
  wire  _T_705 = _T_95 ? 1'h0 : _T_704; // @[Lookup.scala 33:37]
  wire  _T_706 = _T_93 ? 1'h0 : _T_705; // @[Lookup.scala 33:37]
  wire  _T_707 = _T_91 ? 1'h0 : _T_706; // @[Lookup.scala 33:37]
  wire  _T_708 = _T_89 ? 1'h0 : _T_707; // @[Lookup.scala 33:37]
  wire  _T_709 = _T_87 ? 1'h0 : _T_708; // @[Lookup.scala 33:37]
  wire  _T_710 = _T_85 ? 1'h0 : _T_709; // @[Lookup.scala 33:37]
  wire  _T_711 = _T_83 ? 1'h0 : _T_710; // @[Lookup.scala 33:37]
  wire  _T_712 = _T_81 ? 1'h0 : _T_711; // @[Lookup.scala 33:37]
  wire  _T_713 = _T_79 ? 1'h0 : _T_712; // @[Lookup.scala 33:37]
  wire  _T_714 = _T_77 ? 1'h0 : _T_713; // @[Lookup.scala 33:37]
  wire  _T_715 = _T_75 ? 1'h0 : _T_714; // @[Lookup.scala 33:37]
  wire  _T_716 = _T_73 ? 1'h0 : _T_715; // @[Lookup.scala 33:37]
  wire  _T_717 = _T_71 ? 1'h0 : _T_716; // @[Lookup.scala 33:37]
  wire  _T_718 = _T_69 ? 1'h0 : _T_717; // @[Lookup.scala 33:37]
  wire  _T_719 = _T_67 ? 1'h0 : _T_718; // @[Lookup.scala 33:37]
  wire  _T_720 = _T_65 ? 1'h0 : _T_719; // @[Lookup.scala 33:37]
  wire  _T_721 = _T_63 ? 1'h0 : _T_720; // @[Lookup.scala 33:37]
  wire  _T_722 = _T_61 ? 1'h0 : _T_721; // @[Lookup.scala 33:37]
  wire  _T_723 = _T_59 ? 1'h0 : _T_722; // @[Lookup.scala 33:37]
  wire  _T_724 = _T_57 ? 1'h0 : _T_723; // @[Lookup.scala 33:37]
  wire  _T_725 = _T_55 ? 1'h0 : _T_724; // @[Lookup.scala 33:37]
  wire  _T_726 = _T_53 ? 1'h0 : _T_725; // @[Lookup.scala 33:37]
  wire  _T_727 = _T_51 ? 1'h0 : _T_726; // @[Lookup.scala 33:37]
  wire  _T_728 = _T_49 ? 1'h0 : _T_727; // @[Lookup.scala 33:37]
  wire  _T_729 = _T_47 ? 1'h0 : _T_728; // @[Lookup.scala 33:37]
  wire  _T_730 = _T_45 ? 1'h0 : _T_729; // @[Lookup.scala 33:37]
  wire  _T_731 = _T_43 ? 1'h0 : _T_730; // @[Lookup.scala 33:37]
  wire  _T_732 = _T_41 ? 1'h0 : _T_731; // @[Lookup.scala 33:37]
  wire  _T_733 = _T_39 ? 1'h0 : _T_732; // @[Lookup.scala 33:37]
  wire  _T_734 = _T_37 ? 1'h0 : _T_733; // @[Lookup.scala 33:37]
  wire  _T_735 = _T_35 ? 1'h0 : _T_734; // @[Lookup.scala 33:37]
  wire  _T_736 = _T_33 ? 1'h0 : _T_735; // @[Lookup.scala 33:37]
  wire  _T_737 = _T_31 ? 1'h0 : _T_736; // @[Lookup.scala 33:37]
  wire  _T_738 = _T_29 ? 1'h0 : _T_737; // @[Lookup.scala 33:37]
  wire  _T_739 = _T_27 ? 1'h0 : _T_738; // @[Lookup.scala 33:37]
  wire  _T_740 = _T_25 ? 1'h0 : _T_739; // @[Lookup.scala 33:37]
  wire  _T_741 = _T_23 ? 1'h0 : _T_740; // @[Lookup.scala 33:37]
  wire  _T_742 = _T_21 ? 1'h0 : _T_741; // @[Lookup.scala 33:37]
  wire  _T_743 = _T_19 ? 1'h0 : _T_742; // @[Lookup.scala 33:37]
  wire  _T_744 = _T_17 ? 1'h0 : _T_743; // @[Lookup.scala 33:37]
  wire  _T_745 = _T_15 ? 1'h0 : _T_744; // @[Lookup.scala 33:37]
  wire  _T_746 = _T_13 ? 1'h0 : _T_745; // @[Lookup.scala 33:37]
  wire  _T_747 = _T_11 ? 1'h0 : _T_746; // @[Lookup.scala 33:37]
  wire  _T_748 = _T_9 ? 1'h0 : _T_747; // @[Lookup.scala 33:37]
  wire  _T_749 = _T_7 ? 1'h0 : _T_748; // @[Lookup.scala 33:37]
  wire  _T_750 = _T_5 ? 1'h0 : _T_749; // @[Lookup.scala 33:37]
  wire  _T_751 = _T_3 ? 1'h0 : _T_750; // @[Lookup.scala 33:37]
  wire [2:0] _T_752 = _T_101 ? 3'h2 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_753 = _T_99 ? 3'h1 : _T_752; // @[Lookup.scala 33:37]
  wire [2:0] _T_754 = _T_97 ? 3'h0 : _T_753; // @[Lookup.scala 33:37]
  wire [2:0] _T_755 = _T_95 ? 3'h0 : _T_754; // @[Lookup.scala 33:37]
  wire [2:0] _T_756 = _T_93 ? 3'h0 : _T_755; // @[Lookup.scala 33:37]
  wire [2:0] _T_757 = _T_91 ? 3'h0 : _T_756; // @[Lookup.scala 33:37]
  wire [2:0] _T_758 = _T_89 ? 3'h0 : _T_757; // @[Lookup.scala 33:37]
  wire [2:0] _T_759 = _T_87 ? 3'h0 : _T_758; // @[Lookup.scala 33:37]
  wire [2:0] _T_760 = _T_85 ? 3'h0 : _T_759; // @[Lookup.scala 33:37]
  wire [2:0] _T_761 = _T_83 ? 3'h0 : _T_760; // @[Lookup.scala 33:37]
  wire [2:0] _T_762 = _T_81 ? 3'h0 : _T_761; // @[Lookup.scala 33:37]
  wire [2:0] _T_763 = _T_79 ? 3'h0 : _T_762; // @[Lookup.scala 33:37]
  wire [2:0] _T_764 = _T_77 ? 3'h0 : _T_763; // @[Lookup.scala 33:37]
  wire [2:0] _T_765 = _T_75 ? 3'h0 : _T_764; // @[Lookup.scala 33:37]
  wire [2:0] _T_766 = _T_73 ? 3'h0 : _T_765; // @[Lookup.scala 33:37]
  wire [2:0] _T_767 = _T_71 ? 3'h0 : _T_766; // @[Lookup.scala 33:37]
  wire [2:0] _T_768 = _T_69 ? 3'h0 : _T_767; // @[Lookup.scala 33:37]
  wire [2:0] _T_769 = _T_67 ? 3'h0 : _T_768; // @[Lookup.scala 33:37]
  wire [2:0] _T_770 = _T_65 ? 3'h0 : _T_769; // @[Lookup.scala 33:37]
  wire [2:0] _T_771 = _T_63 ? 3'h0 : _T_770; // @[Lookup.scala 33:37]
  wire [2:0] _T_772 = _T_61 ? 3'h0 : _T_771; // @[Lookup.scala 33:37]
  wire [2:0] _T_773 = _T_59 ? 3'h0 : _T_772; // @[Lookup.scala 33:37]
  wire [2:0] _T_774 = _T_57 ? 3'h0 : _T_773; // @[Lookup.scala 33:37]
  wire [2:0] _T_775 = _T_55 ? 3'h0 : _T_774; // @[Lookup.scala 33:37]
  wire [2:0] _T_776 = _T_53 ? 3'h0 : _T_775; // @[Lookup.scala 33:37]
  wire [2:0] _T_777 = _T_51 ? 3'h0 : _T_776; // @[Lookup.scala 33:37]
  wire [2:0] _T_778 = _T_49 ? 3'h0 : _T_777; // @[Lookup.scala 33:37]
  wire [2:0] _T_779 = _T_47 ? 3'h0 : _T_778; // @[Lookup.scala 33:37]
  wire [2:0] _T_780 = _T_45 ? 3'h0 : _T_779; // @[Lookup.scala 33:37]
  wire [2:0] _T_781 = _T_43 ? 3'h0 : _T_780; // @[Lookup.scala 33:37]
  wire [2:0] _T_782 = _T_41 ? 3'h0 : _T_781; // @[Lookup.scala 33:37]
  wire [2:0] _T_783 = _T_39 ? 3'h0 : _T_782; // @[Lookup.scala 33:37]
  wire [2:0] _T_784 = _T_37 ? 3'h0 : _T_783; // @[Lookup.scala 33:37]
  wire [2:0] _T_785 = _T_35 ? 3'h0 : _T_784; // @[Lookup.scala 33:37]
  wire [2:0] _T_786 = _T_33 ? 3'h0 : _T_785; // @[Lookup.scala 33:37]
  wire [2:0] _T_787 = _T_31 ? 3'h0 : _T_786; // @[Lookup.scala 33:37]
  wire [2:0] _T_788 = _T_29 ? 3'h0 : _T_787; // @[Lookup.scala 33:37]
  wire [2:0] _T_789 = _T_27 ? 3'h0 : _T_788; // @[Lookup.scala 33:37]
  wire [2:0] _T_790 = _T_25 ? 3'h0 : _T_789; // @[Lookup.scala 33:37]
  wire [2:0] _T_791 = _T_23 ? 3'h0 : _T_790; // @[Lookup.scala 33:37]
  wire [2:0] _T_792 = _T_21 ? 3'h0 : _T_791; // @[Lookup.scala 33:37]
  wire [2:0] _T_793 = _T_19 ? 3'h0 : _T_792; // @[Lookup.scala 33:37]
  wire [2:0] _T_794 = _T_17 ? 3'h0 : _T_793; // @[Lookup.scala 33:37]
  wire [2:0] _T_795 = _T_15 ? 3'h0 : _T_794; // @[Lookup.scala 33:37]
  wire [2:0] _T_796 = _T_13 ? 3'h0 : _T_795; // @[Lookup.scala 33:37]
  wire [2:0] _T_797 = _T_11 ? 3'h0 : _T_796; // @[Lookup.scala 33:37]
  wire [2:0] _T_798 = _T_9 ? 3'h0 : _T_797; // @[Lookup.scala 33:37]
  wire [2:0] _T_799 = _T_7 ? 3'h0 : _T_798; // @[Lookup.scala 33:37]
  wire [2:0] _T_800 = _T_5 ? 3'h0 : _T_799; // @[Lookup.scala 33:37]
  wire [2:0] _T_801 = _T_3 ? 3'h0 : _T_800; // @[Lookup.scala 33:37]
  assign io_pc_sel = _T_1 ? 2'h0 : _T_151; // @[Lookup.scala 33:37]
  assign io_inst_kill = _T_1 ? 1'h0 : _T_451; // @[Lookup.scala 33:37]
  assign io_A_sel = _T_1 ? 1'h0 : _T_201; // @[Lookup.scala 33:37]
  assign io_B_sel = _T_1 ? 1'h0 : _T_251; // @[Lookup.scala 33:37]
  assign io_imm_sel = _T_1 ? 3'h3 : _T_301; // @[Lookup.scala 33:37]
  assign io_alu_op = _T_1 ? 4'hb : _T_351; // @[Lookup.scala 33:37]
  assign io_br_type = _T_1 ? 3'h0 : _T_401; // @[Lookup.scala 33:37]
  assign io_st_type = _T_1 ? 2'h0 : _T_501; // @[Lookup.scala 33:37]
  assign io_ld_type = _T_1 ? 3'h0 : _T_551; // @[Lookup.scala 33:37]
  assign io_wb_sel = _T_1 ? 2'h0 : _T_601; // @[Lookup.scala 33:37]
  assign io_wb_en = _T_1 | (_T_3 | (_T_5 | (_T_7 | _T_648))); // @[Lookup.scala 33:37]
  assign io_csr_cmd = _T_1 ? 3'h0 : _T_701; // @[Lookup.scala 33:37]
  assign io_illegal = _T_1 ? 1'h0 : _T_751; // @[Lookup.scala 33:37]
  assign io_dfc_cmd = _T_1 ? 3'h0 : _T_801; // @[Lookup.scala 33:37]
endmodule
module Core(
  input         clock,
  input         reset,
  output        io_icache_req_valid,
  output [31:0] io_icache_req_bits_addr,
  input         io_icache_resp_valid,
  input  [31:0] io_icache_resp_bits_data,
  output        io_dcache_abort,
  output        io_dcache_req_valid,
  output [31:0] io_dcache_req_bits_addr,
  output [31:0] io_dcache_req_bits_data,
  output [3:0]  io_dcache_req_bits_mask,
  input         io_dcache_resp_valid,
  input  [31:0] io_dcache_resp_bits_data,
  output        io_table_w_data_valid,
  output [31:0] io_table_w_data_bits_listenAddr,
  output [15:0] io_table_w_data_bits_wPid,
  output        io_table_l_data_valid,
  output [31:0] io_table_l_data_bits_listenAddr,
  output        io_table_e_data_ready,
  input         io_table_e_data_valid,
  input  [15:0] io_table_e_data_bits_pid,
  input         io_table_f_data_valid,
  input         io_table_f_data_bits_full_sig,
  input         io_rxChannel_valid,
  input  [1:0]  pageFault,
  output        io_vmSwitch,
  output [31:0] io_in,
  output        clearPageFault,
  input  [1:0]  pageFault_0,
  output [31:0] satp
);
  wire  dpath_clock; // @[Core.scala 41:21]
  wire  dpath_reset; // @[Core.scala 41:21]
  wire  dpath_io_icache_req_valid; // @[Core.scala 41:21]
  wire [31:0] dpath_io_icache_req_bits_addr; // @[Core.scala 41:21]
  wire  dpath_io_icache_resp_valid; // @[Core.scala 41:21]
  wire [31:0] dpath_io_icache_resp_bits_data; // @[Core.scala 41:21]
  wire  dpath_io_dcache_abort; // @[Core.scala 41:21]
  wire  dpath_io_dcache_req_valid; // @[Core.scala 41:21]
  wire [31:0] dpath_io_dcache_req_bits_addr; // @[Core.scala 41:21]
  wire [31:0] dpath_io_dcache_req_bits_data; // @[Core.scala 41:21]
  wire [3:0] dpath_io_dcache_req_bits_mask; // @[Core.scala 41:21]
  wire  dpath_io_dcache_resp_valid; // @[Core.scala 41:21]
  wire [31:0] dpath_io_dcache_resp_bits_data; // @[Core.scala 41:21]
  wire [31:0] dpath_io_ctrl_inst; // @[Core.scala 41:21]
  wire [1:0] dpath_io_ctrl_pc_sel; // @[Core.scala 41:21]
  wire  dpath_io_ctrl_inst_kill; // @[Core.scala 41:21]
  wire  dpath_io_ctrl_A_sel; // @[Core.scala 41:21]
  wire  dpath_io_ctrl_B_sel; // @[Core.scala 41:21]
  wire [2:0] dpath_io_ctrl_imm_sel; // @[Core.scala 41:21]
  wire [3:0] dpath_io_ctrl_alu_op; // @[Core.scala 41:21]
  wire [2:0] dpath_io_ctrl_br_type; // @[Core.scala 41:21]
  wire [1:0] dpath_io_ctrl_st_type; // @[Core.scala 41:21]
  wire [2:0] dpath_io_ctrl_ld_type; // @[Core.scala 41:21]
  wire [1:0] dpath_io_ctrl_wb_sel; // @[Core.scala 41:21]
  wire  dpath_io_ctrl_wb_en; // @[Core.scala 41:21]
  wire [2:0] dpath_io_ctrl_csr_cmd; // @[Core.scala 41:21]
  wire  dpath_io_ctrl_illegal; // @[Core.scala 41:21]
  wire [2:0] dpath_io_ctrl_dfc_cmd; // @[Core.scala 41:21]
  wire  dpath_io_table_w_data_valid; // @[Core.scala 41:21]
  wire [31:0] dpath_io_table_w_data_bits_listenAddr; // @[Core.scala 41:21]
  wire [15:0] dpath_io_table_w_data_bits_wPid; // @[Core.scala 41:21]
  wire  dpath_io_table_l_data_valid; // @[Core.scala 41:21]
  wire [31:0] dpath_io_table_l_data_bits_listenAddr; // @[Core.scala 41:21]
  wire  dpath_io_table_e_data_ready; // @[Core.scala 41:21]
  wire  dpath_io_table_e_data_valid; // @[Core.scala 41:21]
  wire [15:0] dpath_io_table_e_data_bits_pid; // @[Core.scala 41:21]
  wire  dpath_io_table_f_data_valid; // @[Core.scala 41:21]
  wire  dpath_io_table_f_data_bits_full_sig; // @[Core.scala 41:21]
  wire  dpath_io_rxChannel_valid; // @[Core.scala 41:21]
  wire [1:0] dpath_pageFault; // @[Core.scala 41:21]
  wire  dpath_io_vmSwitch; // @[Core.scala 41:21]
  wire [31:0] dpath_io_in; // @[Core.scala 41:21]
  wire  dpath_clearPageFault; // @[Core.scala 41:21]
  wire [1:0] dpath_pageFault_0; // @[Core.scala 41:21]
  wire [31:0] dpath_satp; // @[Core.scala 41:21]
  wire [31:0] ctrl_io_inst; // @[Core.scala 42:21]
  wire [1:0] ctrl_io_pc_sel; // @[Core.scala 42:21]
  wire  ctrl_io_inst_kill; // @[Core.scala 42:21]
  wire  ctrl_io_A_sel; // @[Core.scala 42:21]
  wire  ctrl_io_B_sel; // @[Core.scala 42:21]
  wire [2:0] ctrl_io_imm_sel; // @[Core.scala 42:21]
  wire [3:0] ctrl_io_alu_op; // @[Core.scala 42:21]
  wire [2:0] ctrl_io_br_type; // @[Core.scala 42:21]
  wire [1:0] ctrl_io_st_type; // @[Core.scala 42:21]
  wire [2:0] ctrl_io_ld_type; // @[Core.scala 42:21]
  wire [1:0] ctrl_io_wb_sel; // @[Core.scala 42:21]
  wire  ctrl_io_wb_en; // @[Core.scala 42:21]
  wire [2:0] ctrl_io_csr_cmd; // @[Core.scala 42:21]
  wire  ctrl_io_illegal; // @[Core.scala 42:21]
  wire [2:0] ctrl_io_dfc_cmd; // @[Core.scala 42:21]
  Datapath dpath ( // @[Core.scala 41:21]
    .clock(dpath_clock),
    .reset(dpath_reset),
    .io_icache_req_valid(dpath_io_icache_req_valid),
    .io_icache_req_bits_addr(dpath_io_icache_req_bits_addr),
    .io_icache_resp_valid(dpath_io_icache_resp_valid),
    .io_icache_resp_bits_data(dpath_io_icache_resp_bits_data),
    .io_dcache_abort(dpath_io_dcache_abort),
    .io_dcache_req_valid(dpath_io_dcache_req_valid),
    .io_dcache_req_bits_addr(dpath_io_dcache_req_bits_addr),
    .io_dcache_req_bits_data(dpath_io_dcache_req_bits_data),
    .io_dcache_req_bits_mask(dpath_io_dcache_req_bits_mask),
    .io_dcache_resp_valid(dpath_io_dcache_resp_valid),
    .io_dcache_resp_bits_data(dpath_io_dcache_resp_bits_data),
    .io_ctrl_inst(dpath_io_ctrl_inst),
    .io_ctrl_pc_sel(dpath_io_ctrl_pc_sel),
    .io_ctrl_inst_kill(dpath_io_ctrl_inst_kill),
    .io_ctrl_A_sel(dpath_io_ctrl_A_sel),
    .io_ctrl_B_sel(dpath_io_ctrl_B_sel),
    .io_ctrl_imm_sel(dpath_io_ctrl_imm_sel),
    .io_ctrl_alu_op(dpath_io_ctrl_alu_op),
    .io_ctrl_br_type(dpath_io_ctrl_br_type),
    .io_ctrl_st_type(dpath_io_ctrl_st_type),
    .io_ctrl_ld_type(dpath_io_ctrl_ld_type),
    .io_ctrl_wb_sel(dpath_io_ctrl_wb_sel),
    .io_ctrl_wb_en(dpath_io_ctrl_wb_en),
    .io_ctrl_csr_cmd(dpath_io_ctrl_csr_cmd),
    .io_ctrl_illegal(dpath_io_ctrl_illegal),
    .io_ctrl_dfc_cmd(dpath_io_ctrl_dfc_cmd),
    .io_table_w_data_valid(dpath_io_table_w_data_valid),
    .io_table_w_data_bits_listenAddr(dpath_io_table_w_data_bits_listenAddr),
    .io_table_w_data_bits_wPid(dpath_io_table_w_data_bits_wPid),
    .io_table_l_data_valid(dpath_io_table_l_data_valid),
    .io_table_l_data_bits_listenAddr(dpath_io_table_l_data_bits_listenAddr),
    .io_table_e_data_ready(dpath_io_table_e_data_ready),
    .io_table_e_data_valid(dpath_io_table_e_data_valid),
    .io_table_e_data_bits_pid(dpath_io_table_e_data_bits_pid),
    .io_table_f_data_valid(dpath_io_table_f_data_valid),
    .io_table_f_data_bits_full_sig(dpath_io_table_f_data_bits_full_sig),
    .io_rxChannel_valid(dpath_io_rxChannel_valid),
    .pageFault(dpath_pageFault),
    .io_vmSwitch(dpath_io_vmSwitch),
    .io_in(dpath_io_in),
    .clearPageFault(dpath_clearPageFault),
    .pageFault_0(dpath_pageFault_0),
    .satp(dpath_satp)
  );
  Control ctrl ( // @[Core.scala 42:21]
    .io_inst(ctrl_io_inst),
    .io_pc_sel(ctrl_io_pc_sel),
    .io_inst_kill(ctrl_io_inst_kill),
    .io_A_sel(ctrl_io_A_sel),
    .io_B_sel(ctrl_io_B_sel),
    .io_imm_sel(ctrl_io_imm_sel),
    .io_alu_op(ctrl_io_alu_op),
    .io_br_type(ctrl_io_br_type),
    .io_st_type(ctrl_io_st_type),
    .io_ld_type(ctrl_io_ld_type),
    .io_wb_sel(ctrl_io_wb_sel),
    .io_wb_en(ctrl_io_wb_en),
    .io_csr_cmd(ctrl_io_csr_cmd),
    .io_illegal(ctrl_io_illegal),
    .io_dfc_cmd(ctrl_io_dfc_cmd)
  );
  assign io_icache_req_valid = dpath_io_icache_req_valid; // @[Core.scala 45:19]
  assign io_icache_req_bits_addr = dpath_io_icache_req_bits_addr; // @[Core.scala 45:19]
  assign io_dcache_abort = dpath_io_dcache_abort; // @[Core.scala 46:19]
  assign io_dcache_req_valid = dpath_io_dcache_req_valid; // @[Core.scala 46:19]
  assign io_dcache_req_bits_addr = dpath_io_dcache_req_bits_addr; // @[Core.scala 46:19]
  assign io_dcache_req_bits_data = dpath_io_dcache_req_bits_data; // @[Core.scala 46:19]
  assign io_dcache_req_bits_mask = dpath_io_dcache_req_bits_mask; // @[Core.scala 46:19]
  assign io_table_w_data_valid = dpath_io_table_w_data_valid; // @[Core.scala 50:14]
  assign io_table_w_data_bits_listenAddr = dpath_io_table_w_data_bits_listenAddr; // @[Core.scala 50:14]
  assign io_table_w_data_bits_wPid = dpath_io_table_w_data_bits_wPid; // @[Core.scala 50:14]
  assign io_table_l_data_valid = dpath_io_table_l_data_valid; // @[Core.scala 51:14]
  assign io_table_l_data_bits_listenAddr = dpath_io_table_l_data_bits_listenAddr; // @[Core.scala 51:14]
  assign io_table_e_data_ready = dpath_io_table_e_data_ready; // @[Core.scala 52:14]
  assign io_vmSwitch = dpath_io_vmSwitch;
  assign io_in = dpath_io_in;
  assign clearPageFault = dpath_clearPageFault;
  assign satp = dpath_satp;
  assign dpath_clock = clock;
  assign dpath_reset = reset;
  assign dpath_io_icache_resp_valid = io_icache_resp_valid; // @[Core.scala 45:19]
  assign dpath_io_icache_resp_bits_data = io_icache_resp_bits_data; // @[Core.scala 45:19]
  assign dpath_io_dcache_resp_valid = io_dcache_resp_valid; // @[Core.scala 46:19]
  assign dpath_io_dcache_resp_bits_data = io_dcache_resp_bits_data; // @[Core.scala 46:19]
  assign dpath_io_ctrl_pc_sel = ctrl_io_pc_sel; // @[Core.scala 47:17]
  assign dpath_io_ctrl_inst_kill = ctrl_io_inst_kill; // @[Core.scala 47:17]
  assign dpath_io_ctrl_A_sel = ctrl_io_A_sel; // @[Core.scala 47:17]
  assign dpath_io_ctrl_B_sel = ctrl_io_B_sel; // @[Core.scala 47:17]
  assign dpath_io_ctrl_imm_sel = ctrl_io_imm_sel; // @[Core.scala 47:17]
  assign dpath_io_ctrl_alu_op = ctrl_io_alu_op; // @[Core.scala 47:17]
  assign dpath_io_ctrl_br_type = ctrl_io_br_type; // @[Core.scala 47:17]
  assign dpath_io_ctrl_st_type = ctrl_io_st_type; // @[Core.scala 47:17]
  assign dpath_io_ctrl_ld_type = ctrl_io_ld_type; // @[Core.scala 47:17]
  assign dpath_io_ctrl_wb_sel = ctrl_io_wb_sel; // @[Core.scala 47:17]
  assign dpath_io_ctrl_wb_en = ctrl_io_wb_en; // @[Core.scala 47:17]
  assign dpath_io_ctrl_csr_cmd = ctrl_io_csr_cmd; // @[Core.scala 47:17]
  assign dpath_io_ctrl_illegal = ctrl_io_illegal; // @[Core.scala 47:17]
  assign dpath_io_ctrl_dfc_cmd = ctrl_io_dfc_cmd; // @[Core.scala 47:17]
  assign dpath_io_table_e_data_valid = io_table_e_data_valid; // @[Core.scala 52:14]
  assign dpath_io_table_e_data_bits_pid = io_table_e_data_bits_pid; // @[Core.scala 52:14]
  assign dpath_io_table_f_data_valid = io_table_f_data_valid; // @[Core.scala 53:14]
  assign dpath_io_table_f_data_bits_full_sig = io_table_f_data_bits_full_sig; // @[Core.scala 53:14]
  assign dpath_io_rxChannel_valid = io_rxChannel_valid;
  assign dpath_pageFault = pageFault;
  assign dpath_pageFault_0 = pageFault_0;
  assign ctrl_io_inst = dpath_io_ctrl_inst; // @[Core.scala 47:17]
endmodule
module Cache(
  input         clock,
  input         reset,
  input         io_cpu_abort,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [31:0] io_cpu_req_bits_data,
  input  [3:0]  io_cpu_req_bits_mask,
  output        io_cpu_resp_valid,
  output [31:0] io_cpu_resp_bits_data,
  input         io_nasti_aw_ready,
  output        io_nasti_aw_valid,
  output [31:0] io_nasti_aw_bits_addr,
  input         io_nasti_w_ready,
  output        io_nasti_w_valid,
  output [31:0] io_nasti_w_bits_data,
  output        io_nasti_w_bits_last,
  output        io_nasti_b_ready,
  input         io_nasti_b_valid,
  input         io_nasti_ar_ready,
  output        io_nasti_ar_valid,
  output [31:0] io_nasti_ar_bits_addr,
  output        io_nasti_r_ready,
  input         io_nasti_r_valid,
  input  [31:0] io_nasti_r_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
`endif // RANDOMIZE_REG_INIT
  reg [29:0] metaMem_tag [0:0]; // @[Cache.scala 69:24]
  wire [29:0] metaMem_tag_rmeta_data; // @[Cache.scala 69:24]
  wire  metaMem_tag_rmeta_addr; // @[Cache.scala 69:24]
  wire [29:0] metaMem_tag_MPORT_1_data; // @[Cache.scala 69:24]
  wire  metaMem_tag_MPORT_1_addr; // @[Cache.scala 69:24]
  wire  metaMem_tag_MPORT_1_mask; // @[Cache.scala 69:24]
  wire  metaMem_tag_MPORT_1_en; // @[Cache.scala 69:24]
  reg  metaMem_tag_rmeta_en_pipe_0;
  reg [7:0] dataMem_0_0 [0:0]; // @[Cache.scala 70:41]
  wire [7:0] dataMem_0_0_MPORT_data; // @[Cache.scala 70:41]
  wire  dataMem_0_0_MPORT_addr; // @[Cache.scala 70:41]
  wire [7:0] dataMem_0_0_MPORT_2_data; // @[Cache.scala 70:41]
  wire  dataMem_0_0_MPORT_2_addr; // @[Cache.scala 70:41]
  wire  dataMem_0_0_MPORT_2_mask; // @[Cache.scala 70:41]
  wire  dataMem_0_0_MPORT_2_en; // @[Cache.scala 70:41]
  reg  dataMem_0_0_MPORT_en_pipe_0;
  reg [7:0] dataMem_0_1 [0:0]; // @[Cache.scala 70:41]
  wire [7:0] dataMem_0_1_MPORT_data; // @[Cache.scala 70:41]
  wire  dataMem_0_1_MPORT_addr; // @[Cache.scala 70:41]
  wire [7:0] dataMem_0_1_MPORT_2_data; // @[Cache.scala 70:41]
  wire  dataMem_0_1_MPORT_2_addr; // @[Cache.scala 70:41]
  wire  dataMem_0_1_MPORT_2_mask; // @[Cache.scala 70:41]
  wire  dataMem_0_1_MPORT_2_en; // @[Cache.scala 70:41]
  reg  dataMem_0_1_MPORT_en_pipe_0;
  reg [7:0] dataMem_0_2 [0:0]; // @[Cache.scala 70:41]
  wire [7:0] dataMem_0_2_MPORT_data; // @[Cache.scala 70:41]
  wire  dataMem_0_2_MPORT_addr; // @[Cache.scala 70:41]
  wire [7:0] dataMem_0_2_MPORT_2_data; // @[Cache.scala 70:41]
  wire  dataMem_0_2_MPORT_2_addr; // @[Cache.scala 70:41]
  wire  dataMem_0_2_MPORT_2_mask; // @[Cache.scala 70:41]
  wire  dataMem_0_2_MPORT_2_en; // @[Cache.scala 70:41]
  reg  dataMem_0_2_MPORT_en_pipe_0;
  reg [7:0] dataMem_0_3 [0:0]; // @[Cache.scala 70:41]
  wire [7:0] dataMem_0_3_MPORT_data; // @[Cache.scala 70:41]
  wire  dataMem_0_3_MPORT_addr; // @[Cache.scala 70:41]
  wire [7:0] dataMem_0_3_MPORT_2_data; // @[Cache.scala 70:41]
  wire  dataMem_0_3_MPORT_2_addr; // @[Cache.scala 70:41]
  wire  dataMem_0_3_MPORT_2_mask; // @[Cache.scala 70:41]
  wire  dataMem_0_3_MPORT_2_en; // @[Cache.scala 70:41]
  reg  dataMem_0_3_MPORT_en_pipe_0;
  reg [2:0] state; // @[Cache.scala 65:22]
  reg  v; // @[Cache.scala 67:25]
  reg  d; // @[Cache.scala 68:25]
  reg [31:0] addr_reg; // @[Cache.scala 72:21]
  reg [31:0] cpu_data; // @[Cache.scala 73:21]
  reg [3:0] cpu_mask; // @[Cache.scala 74:21]
  wire  read_wrap_out = io_nasti_r_ready & io_nasti_r_valid; // @[Decoupled.scala 40:37]
  wire  write_wrap_out = io_nasti_w_ready & io_nasti_w_valid; // @[Decoupled.scala 40:37]
  wire  is_idle = state == 3'h0; // @[Cache.scala 82:25]
  wire  is_read = state == 3'h1; // @[Cache.scala 83:25]
  wire  is_write = state == 3'h2; // @[Cache.scala 84:25]
  wire  is_alloc = state == 3'h6 & read_wrap_out; // @[Cache.scala 85:38]
  reg  is_alloc_reg; // @[Cache.scala 86:29]
  wire [29:0] tag_reg = addr_reg[31:2]; // @[Cache.scala 96:26]
  wire  hit = v & metaMem_tag_rmeta_data == tag_reg; // @[Cache.scala 106:21]
  wire  _T_3 = hit | is_alloc_reg; // @[Cache.scala 89:30]
  wire  _T_6 = is_write & (hit | is_alloc_reg) & ~io_cpu_abort; // @[Cache.scala 89:47]
  wire  wen = is_write & (hit | is_alloc_reg) & ~io_cpu_abort | is_alloc; // @[Cache.scala 89:64]
  wire  _T_9 = ~wen & (is_idle | is_read); // @[Cache.scala 90:18]
  reg  ren_reg; // @[Cache.scala 91:24]
  wire [31:0] rdata = {dataMem_0_3_MPORT_data,dataMem_0_2_MPORT_data,dataMem_0_1_MPORT_data,dataMem_0_0_MPORT_data}; // @[Cache.scala 101:50]
  reg [31:0] rdata_buf; // @[Reg.scala 15:16]
  wire [31:0] _GEN_5 = ren_reg ? rdata : rdata_buf; // @[Reg.scala 16:19 Reg.scala 16:23 Reg.scala 15:16]
  reg [31:0] refill_buf_0; // @[Cache.scala 103:23]
  wire  _T_18 = |cpu_mask; // @[Cache.scala 112:83]
  wire  _T_22 = ~is_alloc; // @[Cache.scala 123:19]
  wire [6:0] _T_23 = {{3'd0}, cpu_mask}; // @[Cache.scala 123:40]
  wire [7:0] _T_24 = {1'b0,$signed(_T_23)}; // @[Cache.scala 123:66]
  wire [7:0] wmask = ~is_alloc ? $signed(_T_24) : $signed(-8'sh1); // @[Cache.scala 123:18]
  wire [31:0] wdata = _T_22 ? cpu_data : io_nasti_r_bits_data; // @[Cache.scala 124:18]
  wire [1:0] _T_38 = _T_22 ? 2'h1 : 2'h2; // @[Cache.scala 129:18]
  wire [1:0] _GEN_22 = wen ? 2'h1 : {{1'd0}, v}; // @[Cache.scala 127:13 Cache.scala 128:7 Cache.scala 67:25]
  wire [1:0] _GEN_23 = wen ? _T_38 : {{1'd0}, d}; // @[Cache.scala 127:13 Cache.scala 129:7 Cache.scala 68:25]
  wire [31:0] _GEN_82 = {tag_reg, 2'h0}; // @[Cache.scala 143:18]
  wire [32:0] _T_48 = {{1'd0}, _GEN_82}; // @[Cache.scala 143:18]
  wire [31:0] _GEN_83 = {metaMem_tag_rmeta_data, 2'h0}; // @[Cache.scala 151:20]
  wire [32:0] _T_52 = {{1'd0}, _GEN_83}; // @[Cache.scala 151:20]
  wire  is_dirty = v & d; // @[Cache.scala 163:29]
  wire  _T_60 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire [2:0] _T_62 = |io_cpu_req_bits_mask ? 3'h2 : 3'h1; // @[Cache.scala 167:21]
  wire  _T_63 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_42 = io_cpu_req_valid ? _T_62 : 3'h0; // @[Cache.scala 172:32 Cache.scala 173:17 Cache.scala 175:17]
  wire  _T_66 = ~is_dirty; // @[Cache.scala 179:30]
  wire  _T_67 = io_nasti_aw_ready & io_nasti_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_68 = io_nasti_ar_ready & io_nasti_ar_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_43 = _T_68 ? 3'h6 : state; // @[Cache.scala 182:40 Cache.scala 183:17 Cache.scala 65:22]
  wire [2:0] _GEN_44 = _T_67 ? 3'h3 : _GEN_43; // @[Cache.scala 180:34 Cache.scala 181:17]
  wire  _GEN_46 = hit ? 1'h0 : is_dirty; // @[Cache.scala 171:17 Cache.scala 152:21 Cache.scala 178:27]
  wire  _GEN_47 = hit ? 1'h0 : ~is_dirty; // @[Cache.scala 171:17 Cache.scala 144:21 Cache.scala 179:27]
  wire  _T_69 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_50 = _T_3 | io_cpu_abort ? 3'h0 : _GEN_44; // @[Cache.scala 188:49 Cache.scala 189:15]
  wire  _GEN_51 = _T_3 | io_cpu_abort ? 1'h0 : is_dirty; // @[Cache.scala 188:49 Cache.scala 152:21 Cache.scala 191:27]
  wire  _GEN_52 = _T_3 | io_cpu_abort ? 1'h0 : _T_66; // @[Cache.scala 188:49 Cache.scala 144:21 Cache.scala 192:27]
  wire  _T_75 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_53 = write_wrap_out ? 3'h4 : state; // @[Cache.scala 202:28 Cache.scala 203:15 Cache.scala 65:22]
  wire  _T_76 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_77 = io_nasti_b_ready & io_nasti_b_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_54 = _T_77 ? 3'h5 : state; // @[Cache.scala 208:31 Cache.scala 209:15 Cache.scala 65:22]
  wire  _T_78 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_80 = 3'h6 == state; // @[Conditional.scala 37:30]
  wire [2:0] _T_82 = _T_18 ? 3'h2 : 3'h0; // @[Cache.scala 220:21]
  wire [2:0] _GEN_56 = read_wrap_out ? _T_82 : state; // @[Cache.scala 219:27 Cache.scala 220:15 Cache.scala 65:22]
  wire [2:0] _GEN_57 = _T_80 ? _GEN_56 : state; // @[Conditional.scala 39:67 Cache.scala 65:22]
  wire [2:0] _GEN_59 = _T_78 ? _GEN_43 : _GEN_57; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_61 = _T_76 ? _GEN_54 : _GEN_59; // @[Conditional.scala 39:67]
  wire  _GEN_62 = _T_76 ? 1'h0 : _T_78; // @[Conditional.scala 39:67 Cache.scala 144:21]
  wire [2:0] _GEN_64 = _T_75 ? _GEN_53 : _GEN_61; // @[Conditional.scala 39:67]
  wire  _GEN_65 = _T_75 ? 1'h0 : _T_76; // @[Conditional.scala 39:67 Cache.scala 160:20]
  wire  _GEN_66 = _T_75 ? 1'h0 : _GEN_62; // @[Conditional.scala 39:67 Cache.scala 144:21]
  wire  _GEN_68 = _T_69 & _GEN_51; // @[Conditional.scala 39:67 Cache.scala 152:21]
  wire  _GEN_69 = _T_69 ? _GEN_52 : _GEN_66; // @[Conditional.scala 39:67]
  wire  _GEN_70 = _T_69 ? 1'h0 : _T_75; // @[Conditional.scala 39:67 Cache.scala 158:20]
  wire  _GEN_71 = _T_69 ? 1'h0 : _GEN_65; // @[Conditional.scala 39:67 Cache.scala 160:20]
  wire  _GEN_73 = _T_63 ? _GEN_46 : _GEN_68; // @[Conditional.scala 39:67]
  wire  _GEN_74 = _T_63 ? _GEN_47 : _GEN_69; // @[Conditional.scala 39:67]
  wire  _GEN_75 = _T_63 ? 1'h0 : _GEN_70; // @[Conditional.scala 39:67 Cache.scala 158:20]
  wire  _GEN_76 = _T_63 ? 1'h0 : _GEN_71; // @[Conditional.scala 39:67 Cache.scala 160:20]
  assign metaMem_tag_rmeta_addr = 1'h0;
  assign metaMem_tag_rmeta_data = metaMem_tag[metaMem_tag_rmeta_addr]; // @[Cache.scala 69:24]
  assign metaMem_tag_MPORT_1_data = addr_reg[31:2];
  assign metaMem_tag_MPORT_1_addr = 1'h0;
  assign metaMem_tag_MPORT_1_mask = 1'h1;
  assign metaMem_tag_MPORT_1_en = wen & is_alloc;
  assign dataMem_0_0_MPORT_addr = 1'h0;
  assign dataMem_0_0_MPORT_data = dataMem_0_0[dataMem_0_0_MPORT_addr]; // @[Cache.scala 70:41]
  assign dataMem_0_0_MPORT_2_data = wdata[7:0];
  assign dataMem_0_0_MPORT_2_addr = 1'h0;
  assign dataMem_0_0_MPORT_2_mask = wmask[0];
  assign dataMem_0_0_MPORT_2_en = _T_6 | is_alloc;
  assign dataMem_0_1_MPORT_addr = 1'h0;
  assign dataMem_0_1_MPORT_data = dataMem_0_1[dataMem_0_1_MPORT_addr]; // @[Cache.scala 70:41]
  assign dataMem_0_1_MPORT_2_data = wdata[15:8];
  assign dataMem_0_1_MPORT_2_addr = 1'h0;
  assign dataMem_0_1_MPORT_2_mask = wmask[1];
  assign dataMem_0_1_MPORT_2_en = _T_6 | is_alloc;
  assign dataMem_0_2_MPORT_addr = 1'h0;
  assign dataMem_0_2_MPORT_data = dataMem_0_2[dataMem_0_2_MPORT_addr]; // @[Cache.scala 70:41]
  assign dataMem_0_2_MPORT_2_data = wdata[23:16];
  assign dataMem_0_2_MPORT_2_addr = 1'h0;
  assign dataMem_0_2_MPORT_2_mask = wmask[2];
  assign dataMem_0_2_MPORT_2_en = _T_6 | is_alloc;
  assign dataMem_0_3_MPORT_addr = 1'h0;
  assign dataMem_0_3_MPORT_data = dataMem_0_3[dataMem_0_3_MPORT_addr]; // @[Cache.scala 70:41]
  assign dataMem_0_3_MPORT_2_data = wdata[31:24];
  assign dataMem_0_3_MPORT_2_addr = 1'h0;
  assign dataMem_0_3_MPORT_2_mask = wmask[3];
  assign dataMem_0_3_MPORT_2_en = _T_6 | is_alloc;
  assign io_cpu_resp_valid = is_idle | is_read & hit | is_alloc_reg & ~(|cpu_mask); // @[Cache.scala 112:54]
  assign io_cpu_resp_bits_data = is_alloc_reg ? refill_buf_0 : _GEN_5; // @[Cache.scala 104:17]
  assign io_nasti_aw_valid = _T_60 ? 1'h0 : _GEN_73; // @[Conditional.scala 40:58 Cache.scala 152:21]
  assign io_nasti_aw_bits_addr = _T_52[31:0]; // @[nasti.scala 158:18 nasti.scala 160:13]
  assign io_nasti_w_valid = _T_60 ? 1'h0 : _GEN_75; // @[Conditional.scala 40:58 Cache.scala 158:20]
  assign io_nasti_w_bits_data = is_alloc_reg ? refill_buf_0 : _GEN_5; // @[Cache.scala 104:17]
  assign io_nasti_w_bits_last = io_nasti_w_ready & io_nasti_w_valid; // @[Decoupled.scala 40:37]
  assign io_nasti_b_ready = _T_60 ? 1'h0 : _GEN_76; // @[Conditional.scala 40:58 Cache.scala 160:20]
  assign io_nasti_ar_valid = _T_60 ? 1'h0 : _GEN_74; // @[Conditional.scala 40:58 Cache.scala 144:21]
  assign io_nasti_ar_bits_addr = _T_48[31:0]; // @[nasti.scala 178:18 nasti.scala 180:13]
  assign io_nasti_r_ready = state == 3'h6; // @[Cache.scala 146:29]
  always @(posedge clock) begin
    if(metaMem_tag_MPORT_1_en & metaMem_tag_MPORT_1_mask) begin
      metaMem_tag[metaMem_tag_MPORT_1_addr] <= metaMem_tag_MPORT_1_data; // @[Cache.scala 69:24]
    end
    metaMem_tag_rmeta_en_pipe_0 <= _T_9 & io_cpu_req_valid;
    if(dataMem_0_0_MPORT_2_en & dataMem_0_0_MPORT_2_mask) begin
      dataMem_0_0[dataMem_0_0_MPORT_2_addr] <= dataMem_0_0_MPORT_2_data; // @[Cache.scala 70:41]
    end
    dataMem_0_0_MPORT_en_pipe_0 <= _T_9 & io_cpu_req_valid;
    if(dataMem_0_1_MPORT_2_en & dataMem_0_1_MPORT_2_mask) begin
      dataMem_0_1[dataMem_0_1_MPORT_2_addr] <= dataMem_0_1_MPORT_2_data; // @[Cache.scala 70:41]
    end
    dataMem_0_1_MPORT_en_pipe_0 <= _T_9 & io_cpu_req_valid;
    if(dataMem_0_2_MPORT_2_en & dataMem_0_2_MPORT_2_mask) begin
      dataMem_0_2[dataMem_0_2_MPORT_2_addr] <= dataMem_0_2_MPORT_2_data; // @[Cache.scala 70:41]
    end
    dataMem_0_2_MPORT_en_pipe_0 <= _T_9 & io_cpu_req_valid;
    if(dataMem_0_3_MPORT_2_en & dataMem_0_3_MPORT_2_mask) begin
      dataMem_0_3[dataMem_0_3_MPORT_2_addr] <= dataMem_0_3_MPORT_2_data; // @[Cache.scala 70:41]
    end
    dataMem_0_3_MPORT_en_pipe_0 <= _T_9 & io_cpu_req_valid;
    if (reset) begin // @[Cache.scala 65:22]
      state <= 3'h0; // @[Cache.scala 65:22]
    end else if (_T_60) begin // @[Conditional.scala 40:58]
      if (io_cpu_req_valid) begin // @[Cache.scala 166:30]
        if (|io_cpu_req_bits_mask) begin // @[Cache.scala 167:21]
          state <= 3'h2;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (_T_63) begin // @[Conditional.scala 39:67]
      if (hit) begin // @[Cache.scala 171:17]
        state <= _GEN_42;
      end else begin
        state <= _GEN_44;
      end
    end else if (_T_69) begin // @[Conditional.scala 39:67]
      state <= _GEN_50;
    end else begin
      state <= _GEN_64;
    end
    if (reset) begin // @[Cache.scala 67:25]
      v <= 1'h0; // @[Cache.scala 67:25]
    end else begin
      v <= _GEN_22[0];
    end
    if (reset) begin // @[Cache.scala 68:25]
      d <= 1'h0; // @[Cache.scala 68:25]
    end else begin
      d <= _GEN_23[0];
    end
    if (io_cpu_resp_valid) begin // @[Cache.scala 114:27]
      addr_reg <= io_cpu_req_bits_addr; // @[Cache.scala 115:15]
    end
    if (io_cpu_resp_valid) begin // @[Cache.scala 114:27]
      cpu_data <= io_cpu_req_bits_data; // @[Cache.scala 116:15]
    end
    if (io_cpu_resp_valid) begin // @[Cache.scala 114:27]
      cpu_mask <= io_cpu_req_bits_mask; // @[Cache.scala 117:15]
    end
    is_alloc_reg <= state == 3'h6 & read_wrap_out; // @[Cache.scala 85:38]
    ren_reg <= ~wen & (is_idle | is_read) & io_cpu_req_valid; // @[Cache.scala 90:42]
    if (ren_reg) begin // @[Reg.scala 16:19]
      rdata_buf <= rdata; // @[Reg.scala 16:23]
    end
    if (read_wrap_out) begin // @[Cache.scala 147:27]
      refill_buf_0 <= io_nasti_r_bits_data; // @[Cache.scala 147:52]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    metaMem_tag[initvar] = _RAND_0[29:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    dataMem_0_0[initvar] = _RAND_2[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    dataMem_0_1[initvar] = _RAND_4[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    dataMem_0_2[initvar] = _RAND_6[7:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    dataMem_0_3[initvar] = _RAND_8[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  metaMem_tag_rmeta_en_pipe_0 = _RAND_1[0:0];
  _RAND_3 = {1{`RANDOM}};
  dataMem_0_0_MPORT_en_pipe_0 = _RAND_3[0:0];
  _RAND_5 = {1{`RANDOM}};
  dataMem_0_1_MPORT_en_pipe_0 = _RAND_5[0:0];
  _RAND_7 = {1{`RANDOM}};
  dataMem_0_2_MPORT_en_pipe_0 = _RAND_7[0:0];
  _RAND_9 = {1{`RANDOM}};
  dataMem_0_3_MPORT_en_pipe_0 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  v = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  d = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  addr_reg = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  cpu_data = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  cpu_mask = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  is_alloc_reg = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ren_reg = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  rdata_buf = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  refill_buf_0 = _RAND_19[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MemArbiter(
  input         clock,
  input         reset,
  output        io_icache_ar_ready,
  input         io_icache_ar_valid,
  input  [31:0] io_icache_ar_bits_addr,
  input         io_icache_r_ready,
  output        io_icache_r_valid,
  output [31:0] io_icache_r_bits_data,
  output        io_dcache_aw_ready,
  input         io_dcache_aw_valid,
  input  [31:0] io_dcache_aw_bits_addr,
  output        io_dcache_w_ready,
  input         io_dcache_w_valid,
  input  [31:0] io_dcache_w_bits_data,
  input         io_dcache_w_bits_last,
  input         io_dcache_b_ready,
  output        io_dcache_b_valid,
  output        io_dcache_ar_ready,
  input         io_dcache_ar_valid,
  input  [31:0] io_dcache_ar_bits_addr,
  input         io_dcache_r_ready,
  output        io_dcache_r_valid,
  output [31:0] io_dcache_r_bits_data,
  input         io_nasti_aw_ready,
  output        io_nasti_aw_valid,
  output [31:0] io_nasti_aw_bits_addr,
  input         io_nasti_w_ready,
  output        io_nasti_w_valid,
  output [31:0] io_nasti_w_bits_data,
  output        io_nasti_w_bits_last,
  output        io_nasti_b_ready,
  input         io_nasti_b_valid,
  input         io_nasti_ar_ready,
  output        io_nasti_ar_valid,
  output [31:0] io_nasti_ar_bits_addr,
  output        io_nasti_r_ready,
  input         io_nasti_r_valid,
  input  [31:0] io_nasti_r_bits_data,
  input         io_nasti_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Tile.scala 22:22]
  wire  _T = state == 3'h0; // @[Tile.scala 27:52]
  wire  _T_4 = state == 3'h3; // @[Tile.scala 33:50]
  wire  _T_8 = state == 3'h4; // @[Tile.scala 39:50]
  wire  _T_18 = ~io_nasti_aw_valid; // @[Tile.scala 51:5]
  wire  _T_19 = (io_icache_ar_valid | io_dcache_ar_valid) & _T_18; // @[Tile.scala 50:67]
  wire  _T_28 = state == 3'h1; // @[Tile.scala 58:50]
  wire  _T_30 = state == 3'h2; // @[Tile.scala 59:50]
  wire  _T_35 = io_dcache_r_ready & _T_30; // @[Tile.scala 61:23]
  wire  _T_37 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_38 = io_dcache_aw_ready & io_dcache_aw_valid; // @[Decoupled.scala 40:37]
  wire  _T_39 = io_dcache_ar_ready & io_dcache_ar_valid; // @[Decoupled.scala 40:37]
  wire  _T_40 = io_icache_ar_ready & io_icache_ar_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_0 = _T_40 ? 3'h1 : state; // @[Tile.scala 70:39 Tile.scala 71:15 Tile.scala 22:22]
  wire  _T_41 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_42 = io_nasti_r_ready & io_nasti_r_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_3 = _T_42 & io_nasti_r_bits_last ? 3'h0 : state; // @[Tile.scala 75:55 Tile.scala 76:15 Tile.scala 22:22]
  wire  _T_44 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_47 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_48 = io_dcache_w_ready & io_dcache_w_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_5 = _T_48 & io_dcache_w_bits_last ? 3'h4 : state; // @[Tile.scala 85:57 Tile.scala 86:15 Tile.scala 22:22]
  wire  _T_50 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_51 = io_nasti_b_ready & io_nasti_b_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_6 = _T_51 ? 3'h0 : state; // @[Tile.scala 90:31 Tile.scala 91:15 Tile.scala 22:22]
  wire [2:0] _GEN_7 = _T_50 ? _GEN_6 : state; // @[Conditional.scala 39:67 Tile.scala 22:22]
  wire [2:0] _GEN_8 = _T_47 ? _GEN_5 : _GEN_7; // @[Conditional.scala 39:67]
  assign io_icache_ar_ready = io_dcache_ar_ready & ~io_dcache_ar_valid; // @[Tile.scala 53:44]
  assign io_icache_r_valid = io_nasti_r_valid & state == 3'h1; // @[Tile.scala 58:41]
  assign io_icache_r_bits_data = io_nasti_r_bits_data; // @[Tile.scala 56:20]
  assign io_dcache_aw_ready = io_nasti_aw_ready & _T; // @[Tile.scala 28:43]
  assign io_dcache_w_ready = io_nasti_w_ready & _T_4; // @[Tile.scala 34:41]
  assign io_dcache_b_valid = io_nasti_b_valid & state == 3'h4; // @[Tile.scala 39:41]
  assign io_dcache_ar_ready = io_nasti_ar_ready & _T_18 & _T; // @[Tile.scala 52:65]
  assign io_dcache_r_valid = io_nasti_r_valid & state == 3'h2; // @[Tile.scala 59:41]
  assign io_dcache_r_bits_data = io_nasti_r_bits_data; // @[Tile.scala 57:20]
  assign io_nasti_aw_valid = io_dcache_aw_valid & state == 3'h0; // @[Tile.scala 27:43]
  assign io_nasti_aw_bits_addr = io_dcache_aw_bits_addr; // @[Tile.scala 26:20]
  assign io_nasti_w_valid = io_dcache_w_valid & state == 3'h3; // @[Tile.scala 33:41]
  assign io_nasti_w_bits_data = io_dcache_w_bits_data; // @[Tile.scala 32:19]
  assign io_nasti_w_bits_last = io_dcache_w_bits_last; // @[Tile.scala 32:19]
  assign io_nasti_b_ready = io_dcache_b_ready & _T_8; // @[Tile.scala 40:41]
  assign io_nasti_ar_valid = _T_19 & _T; // @[Tile.scala 51:24]
  assign io_nasti_ar_bits_addr = io_dcache_ar_valid ? io_dcache_ar_bits_addr : io_icache_ar_bits_addr; // @[Tile.scala 47:8]
  assign io_nasti_r_ready = io_icache_r_ready & _T_28 | _T_35; // @[Tile.scala 60:68]
  always @(posedge clock) begin
    if (reset) begin // @[Tile.scala 22:22]
      state <= 3'h0; // @[Tile.scala 22:22]
    end else if (_T_37) begin // @[Conditional.scala 40:58]
      if (_T_38) begin // @[Tile.scala 66:33]
        state <= 3'h3; // @[Tile.scala 67:15]
      end else if (_T_39) begin // @[Tile.scala 68:39]
        state <= 3'h2; // @[Tile.scala 69:15]
      end else begin
        state <= _GEN_0;
      end
    end else if (_T_41) begin // @[Conditional.scala 39:67]
      state <= _GEN_3;
    end else if (_T_44) begin // @[Conditional.scala 39:67]
      state <= _GEN_3;
    end else begin
      state <= _GEN_8;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Selector(
  input         clock,
  input         reset,
  input         io_cpu_abort,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [31:0] io_cpu_req_bits_data,
  input  [3:0]  io_cpu_req_bits_mask,
  output        io_cpu_resp_valid,
  output [31:0] io_cpu_resp_bits_data,
  output        io_dcache_abort,
  output        io_dcache_req_valid,
  output [31:0] io_dcache_req_bits_addr,
  output [31:0] io_dcache_req_bits_data,
  output [3:0]  io_dcache_req_bits_mask,
  input         io_dcache_resp_valid,
  input  [31:0] io_dcache_resp_bits_data,
  output        io_devices_req_valid,
  output [31:0] io_devices_req_bits_addr,
  output [31:0] io_devices_req_bits_data,
  output [3:0]  io_devices_req_bits_mask,
  input         io_devices_resp_valid,
  input  [31:0] io_devices_resp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] addr; // @[Selector.scala 22:21]
  wire [31:0] _T = io_cpu_req_bits_addr & 32'hf0000000; // @[Selector.scala 32:48]
  wire  _T_1 = 32'h10000000 == _T; // @[Selector.scala 32:48]
  wire [31:0] _T_7 = addr & 32'hf0000000; // @[Selector.scala 41:11]
  wire  _T_8 = 32'h10000000 == _T_7; // @[Selector.scala 41:11]
  assign io_cpu_resp_valid = _T_8 ? io_devices_resp_valid : io_dcache_resp_valid; // @[Mux.scala 98:16]
  assign io_cpu_resp_bits_data = _T_8 ? io_devices_resp_bits_data : io_dcache_resp_bits_data; // @[Mux.scala 98:16]
  assign io_dcache_abort = io_cpu_abort; // @[Selector.scala 47:19]
  assign io_dcache_req_valid = ~(32'h10000000 == _T) & io_cpu_req_valid; // @[Selector.scala 32:70]
  assign io_dcache_req_bits_addr = io_cpu_req_bits_addr; // @[Selector.scala 29:27]
  assign io_dcache_req_bits_data = io_cpu_req_bits_data; // @[Selector.scala 30:27]
  assign io_dcache_req_bits_mask = io_cpu_req_bits_mask; // @[Selector.scala 31:27]
  assign io_devices_req_valid = _T_1 & io_cpu_req_valid; // @[Selector.scala 38:71]
  assign io_devices_req_bits_addr = io_cpu_req_bits_addr; // @[Selector.scala 35:28]
  assign io_devices_req_bits_data = io_cpu_req_bits_data; // @[Selector.scala 36:28]
  assign io_devices_req_bits_mask = io_cpu_req_bits_mask; // @[Selector.scala 37:28]
  always @(posedge clock) begin
    if (reset) begin // @[Selector.scala 22:21]
      addr <= 32'h0; // @[Selector.scala 22:21]
    end else if (io_cpu_req_valid) begin // @[Selector.scala 24:27]
      addr <= io_cpu_req_bits_addr; // @[Selector.scala 25:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MMU(
  input         clock,
  input         reset,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  output        io_cpu_resp_valid,
  output [31:0] io_cpu_resp_bits_data,
  output        io_cache_req_valid,
  output [31:0] io_cache_req_bits_addr,
  input         io_cache_resp_valid,
  input  [31:0] io_cache_resp_bits_data,
  input         vmSwitch_0,
  input  [31:0] csrWdata_0,
  input         clearPageFault_0,
  output [1:0]  pageFault_1,
  input  [31:0] satp_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] satp = vmSwitch_0 ? csrWdata_0 : satp_0; // @[MMU.scala 32:17]
  reg [31:0] rdata; // @[MMU.scala 36:22]
  wire  MODE = satp[31]; // @[MMU.scala 39:18]
  wire [21:0] PPN = satp[21:0]; // @[MMU.scala 41:17]
  reg [31:0] cpu_addr; // @[Reg.scala 15:16]
  wire [9:0] VPN1 = cpu_addr[31:22]; // @[MMU.scala 45:28]
  wire [9:0] VPN0 = cpu_addr[21:12]; // @[MMU.scala 46:28]
  wire [11:0] pageOffest = cpu_addr[11:0]; // @[MMU.scala 47:28]
  wire [11:0] PPN1 = rdata[31:20]; // @[MMU.scala 50:19]
  wire [9:0] PPN0 = rdata[19:10]; // @[MMU.scala 51:19]
  wire  V = rdata[0]; // @[MMU.scala 65:16]
  wire [34:0] _T = PPN * 13'h1000; // @[MMU.scala 70:32]
  wire [12:0] _T_1 = VPN1 * 3'h4; // @[MMU.scala 70:50]
  wire [34:0] _GEN_87 = {{22'd0}, _T_1}; // @[MMU.scala 70:43]
  wire [34:0] LevelOnePTEAddress = _T + _GEN_87; // @[MMU.scala 70:43]
  wire [21:0] _T_3 = {PPN1,PPN0}; // @[Cat.scala 30:58]
  wire [34:0] _T_4 = _T_3 * 13'h1000; // @[MMU.scala 71:44]
  wire [12:0] _T_5 = VPN0 * 3'h4; // @[MMU.scala 71:62]
  wire [34:0] _GEN_88 = {{22'd0}, _T_5}; // @[MMU.scala 71:55]
  wire [34:0] LevelTwoPTEAddress = _T_4 + _GEN_88; // @[MMU.scala 71:55]
  reg [3:0] state; // @[MMU.scala 75:22]
  reg [31:0] cacheReqAddr; // @[MMU.scala 78:29]
  wire  _T_7 = ~MODE; // @[MMU.scala 83:38]
  wire [31:0] _T_8 = ~MODE ? io_cpu_req_bits_addr : cacheReqAddr; // @[MMU.scala 83:32]
  reg [1:0] pageFault; // @[MMU.scala 97:26]
  wire [33:0] physicalAddress = {PPN1,PPN0,pageOffest}; // @[Cat.scala 30:58]
  reg [31:0] cpuRespData; // @[MMU.scala 108:28]
  wire  _T_27 = 4'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_32 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_33 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_6 = io_cache_resp_valid ? io_cache_resp_bits_data : rdata; // @[MMU.scala 131:32 MMU.scala 132:15 MMU.scala 36:22]
  wire [3:0] _GEN_7 = io_cache_resp_valid ? 4'h3 : state; // @[MMU.scala 131:32 MMU.scala 133:15 MMU.scala 75:22]
  wire  _T_34 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire [34:0] _GEN_8 = V ? LevelTwoPTEAddress : {{3'd0}, _T_8}; // @[MMU.scala 140:31 MMU.scala 141:34 MMU.scala 83:26]
  wire  _GEN_9 = V | _T_7 & io_cpu_req_valid; // @[MMU.scala 140:31 MMU.scala 142:30 MMU.scala 87:22]
  wire [3:0] _GEN_10 = V ? 4'h4 : 4'h0; // @[MMU.scala 140:31 MMU.scala 143:17 MMU.scala 150:15]
  wire [1:0] _GEN_11 = V ? pageFault : 2'h1; // @[MMU.scala 140:31 MMU.scala 97:26 MMU.scala 147:19]
  wire  _T_39 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_16 = io_cache_resp_valid ? 4'h5 : state; // @[MMU.scala 154:32 MMU.scala 156:15 MMU.scala 75:22]
  wire  _T_40 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire [33:0] _GEN_17 = V ? physicalAddress : {{2'd0}, _T_8}; // @[MMU.scala 163:31 MMU.scala 166:34 MMU.scala 83:26]
  wire [3:0] _GEN_21 = V ? 4'h7 : 4'h0; // @[MMU.scala 163:31 MMU.scala 171:17 MMU.scala 179:17]
  wire  _T_47 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_29 = io_cache_resp_valid ? 4'h0 : state; // @[MMU.scala 187:37 MMU.scala 188:19 MMU.scala 75:22]
  wire  _T_48 = 4'h7 == state; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_31 = io_cache_resp_valid ? io_cache_resp_bits_data : cpuRespData; // @[MMU.scala 197:37 MMU.scala 198:25 MMU.scala 108:28]
  wire [3:0] _GEN_33 = _T_48 ? _GEN_29 : state; // @[Conditional.scala 39:67 MMU.scala 75:22]
  wire [31:0] _GEN_34 = _T_48 ? _GEN_31 : cpuRespData; // @[Conditional.scala 39:67 MMU.scala 108:28]
  wire [3:0] _GEN_35 = _T_47 ? _GEN_29 : _GEN_33; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_36 = _T_47 ? cpuRespData : _GEN_34; // @[Conditional.scala 39:67 MMU.scala 108:28]
  wire [3:0] _GEN_37 = _T_40 ? _GEN_21 : _GEN_35; // @[Conditional.scala 39:67]
  wire [33:0] _GEN_38 = _T_40 ? _GEN_17 : {{2'd0}, _T_8}; // @[Conditional.scala 39:67 MMU.scala 83:26]
  wire  _GEN_41 = _T_40 ? _GEN_9 : _T_7 & io_cpu_req_valid; // @[Conditional.scala 39:67 MMU.scala 87:22]
  wire [1:0] _GEN_42 = _T_40 ? _GEN_11 : pageFault; // @[Conditional.scala 39:67 MMU.scala 97:26]
  wire [31:0] _GEN_43 = _T_40 ? cpuRespData : _GEN_36; // @[Conditional.scala 39:67 MMU.scala 108:28]
  wire [31:0] _GEN_44 = _T_39 ? _GEN_6 : rdata; // @[Conditional.scala 39:67 MMU.scala 36:22]
  wire [3:0] _GEN_45 = _T_39 ? _GEN_16 : _GEN_37; // @[Conditional.scala 39:67]
  wire [33:0] _GEN_46 = _T_39 ? {{2'd0}, _T_8} : _GEN_38; // @[Conditional.scala 39:67 MMU.scala 83:26]
  wire  _GEN_49 = _T_39 ? _T_7 & io_cpu_req_valid : _GEN_41; // @[Conditional.scala 39:67 MMU.scala 87:22]
  wire [1:0] _GEN_50 = _T_39 ? pageFault : _GEN_42; // @[Conditional.scala 39:67 MMU.scala 97:26]
  wire [31:0] _GEN_51 = _T_39 ? cpuRespData : _GEN_43; // @[Conditional.scala 39:67 MMU.scala 108:28]
  wire [3:0] _GEN_52 = _T_34 ? _GEN_10 : _GEN_45; // @[Conditional.scala 39:67]
  wire [34:0] _GEN_53 = _T_34 ? _GEN_8 : {{1'd0}, _GEN_46}; // @[Conditional.scala 39:67]
  wire  _GEN_54 = _T_34 ? _GEN_9 : _GEN_49; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_55 = _T_34 ? _GEN_11 : _GEN_50; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_56 = _T_34 ? rdata : _GEN_44; // @[Conditional.scala 39:67 MMU.scala 36:22]
  wire [31:0] _GEN_59 = _T_34 ? cpuRespData : _GEN_51; // @[Conditional.scala 39:67 MMU.scala 108:28]
  wire [34:0] _GEN_62 = _T_33 ? {{3'd0}, _T_8} : _GEN_53; // @[Conditional.scala 39:67 MMU.scala 83:26]
  wire  _GEN_63 = _T_33 ? _T_7 & io_cpu_req_valid : _GEN_54; // @[Conditional.scala 39:67 MMU.scala 87:22]
  wire [34:0] _GEN_68 = _T_32 ? LevelOnePTEAddress : _GEN_62; // @[Conditional.scala 39:67 MMU.scala 126:30]
  wire  _GEN_69 = _T_32 | _GEN_63; // @[Conditional.scala 39:67 MMU.scala 127:26]
  wire [34:0] _GEN_81 = _T_27 ? {{3'd0}, _T_8} : _GEN_68; // @[Conditional.scala 40:58 MMU.scala 83:26]
  assign io_cpu_resp_valid = _T_7 ? io_cache_resp_valid : state == 4'h0; // @[MMU.scala 110:27]
  assign io_cpu_resp_bits_data = _T_7 ? io_cache_resp_bits_data : cpuRespData; // @[MMU.scala 109:31]
  assign io_cache_req_valid = _T_27 ? _T_7 & io_cpu_req_valid : _GEN_69; // @[Conditional.scala 40:58 MMU.scala 87:22]
  assign io_cache_req_bits_addr = _GEN_81[31:0];
  assign pageFault_1 = pageFault;
  always @(posedge clock) begin
    if (reset) begin // @[MMU.scala 36:22]
      rdata <= 32'h0; // @[MMU.scala 36:22]
    end else if (!(_T_27)) begin // @[Conditional.scala 40:58]
      if (!(_T_32)) begin // @[Conditional.scala 39:67]
        if (_T_33) begin // @[Conditional.scala 39:67]
          rdata <= _GEN_6;
        end else begin
          rdata <= _GEN_56;
        end
      end
    end
    if (io_cpu_req_valid) begin // @[Reg.scala 16:19]
      cpu_addr <= io_cpu_req_bits_addr; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[MMU.scala 75:22]
      state <= 4'h0; // @[MMU.scala 75:22]
    end else if (_T_27) begin // @[Conditional.scala 40:58]
      if (io_cpu_req_valid & MODE) begin // @[MMU.scala 116:62]
        state <= 4'h1; // @[MMU.scala 121:15]
      end
    end else if (_T_32) begin // @[Conditional.scala 39:67]
      state <= 4'h2; // @[MMU.scala 128:13]
    end else if (_T_33) begin // @[Conditional.scala 39:67]
      state <= _GEN_7;
    end else begin
      state <= _GEN_52;
    end
    if (reset) begin // @[MMU.scala 78:29]
      cacheReqAddr <= 32'h0; // @[MMU.scala 78:29]
    end else if (_T_27) begin // @[Conditional.scala 40:58]
      if (io_cpu_req_valid & MODE) begin // @[MMU.scala 116:62]
        cacheReqAddr <= io_cpu_req_bits_addr; // @[MMU.scala 118:22]
      end
    end
    if (reset) begin // @[MMU.scala 97:26]
      pageFault <= 2'h0; // @[MMU.scala 97:26]
    end else if (_T_27) begin // @[Conditional.scala 40:58]
      if (clearPageFault_0) begin // @[MMU.scala 115:27]
        pageFault <= 2'h0; // @[MMU.scala 115:38]
      end
    end else if (!(_T_32)) begin // @[Conditional.scala 39:67]
      if (!(_T_33)) begin // @[Conditional.scala 39:67]
        pageFault <= _GEN_55;
      end
    end
    if (reset) begin // @[MMU.scala 108:28]
      cpuRespData <= 32'h0; // @[MMU.scala 108:28]
    end else if (!(_T_27)) begin // @[Conditional.scala 40:58]
      if (!(_T_32)) begin // @[Conditional.scala 39:67]
        if (!(_T_33)) begin // @[Conditional.scala 39:67]
          cpuRespData <= _GEN_59;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rdata = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cpu_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  cacheReqAddr = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  pageFault = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  cpuRespData = _RAND_5[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MMU_1(
  input         clock,
  input         reset,
  input         io_cpu_abort,
  input         io_cpu_req_valid,
  input  [31:0] io_cpu_req_bits_addr,
  input  [31:0] io_cpu_req_bits_data,
  input  [3:0]  io_cpu_req_bits_mask,
  output        io_cpu_resp_valid,
  output [31:0] io_cpu_resp_bits_data,
  output        io_cache_abort,
  output        io_cache_req_valid,
  output [31:0] io_cache_req_bits_addr,
  output [31:0] io_cache_req_bits_data,
  output [3:0]  io_cache_req_bits_mask,
  input         io_cache_resp_valid,
  input  [31:0] io_cache_resp_bits_data,
  output [1:0]  pageFault_0,
  input         vmSwitch_0,
  input  [31:0] csrWdata_0,
  input         clearPageFault_0,
  input  [31:0] satp_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] satp = vmSwitch_0 ? csrWdata_0 : satp_0; // @[MMU.scala 32:17]
  reg [31:0] rdata; // @[MMU.scala 36:22]
  wire  MODE = satp[31]; // @[MMU.scala 39:18]
  wire [21:0] PPN = satp[21:0]; // @[MMU.scala 41:17]
  reg [31:0] cpu_addr; // @[Reg.scala 15:16]
  wire [9:0] VPN1 = cpu_addr[31:22]; // @[MMU.scala 45:28]
  wire [9:0] VPN0 = cpu_addr[21:12]; // @[MMU.scala 46:28]
  wire [11:0] pageOffest = cpu_addr[11:0]; // @[MMU.scala 47:28]
  wire [11:0] PPN1 = rdata[31:20]; // @[MMU.scala 50:19]
  wire [9:0] PPN0 = rdata[19:10]; // @[MMU.scala 51:19]
  wire  V = rdata[0]; // @[MMU.scala 65:16]
  wire [34:0] _T = PPN * 13'h1000; // @[MMU.scala 70:32]
  wire [12:0] _T_1 = VPN1 * 3'h4; // @[MMU.scala 70:50]
  wire [34:0] _GEN_87 = {{22'd0}, _T_1}; // @[MMU.scala 70:43]
  wire [34:0] LevelOnePTEAddress = _T + _GEN_87; // @[MMU.scala 70:43]
  wire [21:0] _T_3 = {PPN1,PPN0}; // @[Cat.scala 30:58]
  wire [34:0] _T_4 = _T_3 * 13'h1000; // @[MMU.scala 71:44]
  wire [12:0] _T_5 = VPN0 * 3'h4; // @[MMU.scala 71:62]
  wire [34:0] _GEN_88 = {{22'd0}, _T_5}; // @[MMU.scala 71:55]
  wire [34:0] LevelTwoPTEAddress = _T_4 + _GEN_88; // @[MMU.scala 71:55]
  reg [3:0] state; // @[MMU.scala 75:22]
  reg [31:0] cacheReqAddr; // @[MMU.scala 78:29]
  reg [31:0] cacheReqData; // @[MMU.scala 79:30]
  reg [3:0] cacheReqMask; // @[MMU.scala 80:30]
  wire  _T_7 = ~MODE; // @[MMU.scala 83:38]
  wire [31:0] _T_8 = ~MODE ? io_cpu_req_bits_addr : cacheReqAddr; // @[MMU.scala 83:32]
  wire [31:0] _T_10 = _T_7 ? io_cpu_req_bits_data : cacheReqData; // @[MMU.scala 84:32]
  wire  _T_13 = ~io_cpu_abort; // @[MMU.scala 86:69]
  wire [3:0] _T_15 = state == 4'h5 & ~io_cpu_abort ? io_cpu_req_bits_mask : 4'h0; // @[MMU.scala 86:36]
  wire [3:0] _T_16 = _T_7 ? io_cpu_req_bits_mask : _T_15; // @[MMU.scala 85:32]
  reg [1:0] pageFault; // @[MMU.scala 97:26]
  wire  isLoad = ^io_cpu_req_bits_mask; // @[MMU.scala 99:73]
  wire  isStore = ~isLoad; // @[MMU.scala 100:49]
  wire [33:0] physicalAddress = {PPN1,PPN0,pageOffest}; // @[Cat.scala 30:58]
  reg [31:0] cpuRespData; // @[MMU.scala 108:28]
  wire  _T_27 = 4'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_32 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_33 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_6 = io_cache_resp_valid ? io_cache_resp_bits_data : rdata; // @[MMU.scala 131:32 MMU.scala 132:15 MMU.scala 36:22]
  wire [3:0] _GEN_7 = io_cache_resp_valid ? 4'h3 : state; // @[MMU.scala 131:32 MMU.scala 133:15 MMU.scala 75:22]
  wire  _T_34 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire [1:0] _T_36 = isStore ? 2'h3 : 2'h0; // @[MMU.scala 149:28]
  wire [1:0] _T_37 = isLoad ? 2'h2 : _T_36; // @[MMU.scala 148:28]
  wire [34:0] _GEN_8 = V ? LevelTwoPTEAddress : {{3'd0}, _T_8}; // @[MMU.scala 140:31 MMU.scala 141:34 MMU.scala 83:26]
  wire  _GEN_9 = V | _T_7 & io_cpu_req_valid; // @[MMU.scala 140:31 MMU.scala 142:30 MMU.scala 87:22]
  wire [3:0] _GEN_10 = V ? 4'h4 : 4'h0; // @[MMU.scala 140:31 MMU.scala 143:17 MMU.scala 150:15]
  wire [1:0] _GEN_11 = V ? pageFault : _T_37; // @[MMU.scala 140:31 MMU.scala 97:26 MMU.scala 147:19]
  wire [3:0] _GEN_12 = io_cpu_abort ? 4'h0 : _GEN_10; // @[MMU.scala 137:26 MMU.scala 138:15]
  wire [34:0] _GEN_13 = io_cpu_abort ? {{3'd0}, _T_8} : _GEN_8; // @[MMU.scala 137:26 MMU.scala 83:26]
  wire  _GEN_14 = io_cpu_abort ? _T_7 & io_cpu_req_valid : _GEN_9; // @[MMU.scala 137:26 MMU.scala 87:22]
  wire [1:0] _GEN_15 = io_cpu_abort ? pageFault : _GEN_11; // @[MMU.scala 137:26 MMU.scala 97:26]
  wire  _T_39 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_16 = io_cache_resp_valid ? 4'h5 : state; // @[MMU.scala 154:32 MMU.scala 156:15 MMU.scala 75:22]
  wire  _T_40 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire [3:0] _T_43 = |io_cpu_req_bits_mask ? 4'h6 : 4'h7; // @[MMU.scala 171:23]
  wire [33:0] _GEN_17 = V ? physicalAddress : {{2'd0}, _T_8}; // @[MMU.scala 163:31 MMU.scala 166:34 MMU.scala 83:26]
  wire [31:0] _GEN_18 = V ? cacheReqData : _T_10; // @[MMU.scala 163:31 MMU.scala 167:34 MMU.scala 84:26]
  wire [3:0] _GEN_19 = V ? cacheReqMask : _T_16; // @[MMU.scala 163:31 MMU.scala 168:34 MMU.scala 85:26]
  wire [3:0] _GEN_21 = V ? _T_43 : 4'h0; // @[MMU.scala 163:31 MMU.scala 171:17 MMU.scala 179:17]
  wire [3:0] _GEN_23 = io_cpu_abort ? 4'h0 : _GEN_21; // @[MMU.scala 160:26 MMU.scala 161:15]
  wire [33:0] _GEN_24 = io_cpu_abort ? {{2'd0}, _T_8} : _GEN_17; // @[MMU.scala 160:26 MMU.scala 83:26]
  wire [31:0] _GEN_25 = io_cpu_abort ? _T_10 : _GEN_18; // @[MMU.scala 160:26 MMU.scala 84:26]
  wire [3:0] _GEN_26 = io_cpu_abort ? _T_16 : _GEN_19; // @[MMU.scala 160:26 MMU.scala 85:26]
  wire  _T_47 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_29 = io_cache_resp_valid ? 4'h0 : state; // @[MMU.scala 187:37 MMU.scala 188:19 MMU.scala 75:22]
  wire [3:0] _GEN_30 = io_cpu_abort ? 4'h0 : _GEN_29; // @[MMU.scala 183:26 MMU.scala 184:15]
  wire  _T_48 = 4'h7 == state; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_31 = io_cache_resp_valid ? io_cache_resp_bits_data : cpuRespData; // @[MMU.scala 197:37 MMU.scala 198:25 MMU.scala 108:28]
  wire [31:0] _GEN_32 = io_cpu_abort ? cpuRespData : _GEN_31; // @[MMU.scala 193:26 MMU.scala 108:28]
  wire [3:0] _GEN_33 = _T_48 ? _GEN_30 : state; // @[Conditional.scala 39:67 MMU.scala 75:22]
  wire [31:0] _GEN_34 = _T_48 ? _GEN_32 : cpuRespData; // @[Conditional.scala 39:67 MMU.scala 108:28]
  wire [3:0] _GEN_35 = _T_47 ? _GEN_30 : _GEN_33; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_36 = _T_47 ? cpuRespData : _GEN_34; // @[Conditional.scala 39:67 MMU.scala 108:28]
  wire [3:0] _GEN_37 = _T_40 ? _GEN_23 : _GEN_35; // @[Conditional.scala 39:67]
  wire [33:0] _GEN_38 = _T_40 ? _GEN_24 : {{2'd0}, _T_8}; // @[Conditional.scala 39:67 MMU.scala 83:26]
  wire [31:0] _GEN_39 = _T_40 ? _GEN_25 : _T_10; // @[Conditional.scala 39:67 MMU.scala 84:26]
  wire [3:0] _GEN_40 = _T_40 ? _GEN_26 : _T_16; // @[Conditional.scala 39:67 MMU.scala 85:26]
  wire  _GEN_41 = _T_40 ? _GEN_14 : _T_7 & io_cpu_req_valid; // @[Conditional.scala 39:67 MMU.scala 87:22]
  wire [1:0] _GEN_42 = _T_40 ? _GEN_15 : pageFault; // @[Conditional.scala 39:67 MMU.scala 97:26]
  wire [31:0] _GEN_43 = _T_40 ? cpuRespData : _GEN_36; // @[Conditional.scala 39:67 MMU.scala 108:28]
  wire [31:0] _GEN_44 = _T_39 ? _GEN_6 : rdata; // @[Conditional.scala 39:67 MMU.scala 36:22]
  wire [3:0] _GEN_45 = _T_39 ? _GEN_16 : _GEN_37; // @[Conditional.scala 39:67]
  wire [33:0] _GEN_46 = _T_39 ? {{2'd0}, _T_8} : _GEN_38; // @[Conditional.scala 39:67 MMU.scala 83:26]
  wire [31:0] _GEN_47 = _T_39 ? _T_10 : _GEN_39; // @[Conditional.scala 39:67 MMU.scala 84:26]
  wire [3:0] _GEN_48 = _T_39 ? _T_16 : _GEN_40; // @[Conditional.scala 39:67 MMU.scala 85:26]
  wire  _GEN_49 = _T_39 ? _T_7 & io_cpu_req_valid : _GEN_41; // @[Conditional.scala 39:67 MMU.scala 87:22]
  wire [1:0] _GEN_50 = _T_39 ? pageFault : _GEN_42; // @[Conditional.scala 39:67 MMU.scala 97:26]
  wire [31:0] _GEN_51 = _T_39 ? cpuRespData : _GEN_43; // @[Conditional.scala 39:67 MMU.scala 108:28]
  wire [3:0] _GEN_52 = _T_34 ? _GEN_12 : _GEN_45; // @[Conditional.scala 39:67]
  wire [34:0] _GEN_53 = _T_34 ? _GEN_13 : {{1'd0}, _GEN_46}; // @[Conditional.scala 39:67]
  wire  _GEN_54 = _T_34 ? _GEN_14 : _GEN_49; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_55 = _T_34 ? _GEN_15 : _GEN_50; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_56 = _T_34 ? rdata : _GEN_44; // @[Conditional.scala 39:67 MMU.scala 36:22]
  wire [31:0] _GEN_57 = _T_34 ? _T_10 : _GEN_47; // @[Conditional.scala 39:67 MMU.scala 84:26]
  wire [3:0] _GEN_58 = _T_34 ? _T_16 : _GEN_48; // @[Conditional.scala 39:67 MMU.scala 85:26]
  wire [31:0] _GEN_59 = _T_34 ? cpuRespData : _GEN_51; // @[Conditional.scala 39:67 MMU.scala 108:28]
  wire [34:0] _GEN_62 = _T_33 ? {{3'd0}, _T_8} : _GEN_53; // @[Conditional.scala 39:67 MMU.scala 83:26]
  wire  _GEN_63 = _T_33 ? _T_7 & io_cpu_req_valid : _GEN_54; // @[Conditional.scala 39:67 MMU.scala 87:22]
  wire [31:0] _GEN_65 = _T_33 ? _T_10 : _GEN_57; // @[Conditional.scala 39:67 MMU.scala 84:26]
  wire [3:0] _GEN_66 = _T_33 ? _T_16 : _GEN_58; // @[Conditional.scala 39:67 MMU.scala 85:26]
  wire [34:0] _GEN_68 = _T_32 ? LevelOnePTEAddress : _GEN_62; // @[Conditional.scala 39:67 MMU.scala 126:30]
  wire  _GEN_69 = _T_32 | _GEN_63; // @[Conditional.scala 39:67 MMU.scala 127:26]
  wire [31:0] _GEN_73 = _T_32 ? _T_10 : _GEN_65; // @[Conditional.scala 39:67 MMU.scala 84:26]
  wire [3:0] _GEN_74 = _T_32 ? _T_16 : _GEN_66; // @[Conditional.scala 39:67 MMU.scala 85:26]
  wire [34:0] _GEN_81 = _T_27 ? {{3'd0}, _T_8} : _GEN_68; // @[Conditional.scala 40:58 MMU.scala 83:26]
  assign io_cpu_resp_valid = _T_7 ? io_cache_resp_valid : state == 4'h0; // @[MMU.scala 110:27]
  assign io_cpu_resp_bits_data = _T_7 ? io_cache_resp_bits_data : cpuRespData; // @[MMU.scala 109:31]
  assign io_cache_abort = io_cpu_abort; // @[MMU.scala 88:18]
  assign io_cache_req_valid = _T_27 ? _T_7 & io_cpu_req_valid : _GEN_69; // @[Conditional.scala 40:58 MMU.scala 87:22]
  assign io_cache_req_bits_addr = _GEN_81[31:0];
  assign io_cache_req_bits_data = _T_27 ? _T_10 : _GEN_73; // @[Conditional.scala 40:58 MMU.scala 84:26]
  assign io_cache_req_bits_mask = _T_27 ? _T_16 : _GEN_74; // @[Conditional.scala 40:58 MMU.scala 85:26]
  assign pageFault_0 = pageFault;
  always @(posedge clock) begin
    if (reset) begin // @[MMU.scala 36:22]
      rdata <= 32'h0; // @[MMU.scala 36:22]
    end else if (!(_T_27)) begin // @[Conditional.scala 40:58]
      if (!(_T_32)) begin // @[Conditional.scala 39:67]
        if (_T_33) begin // @[Conditional.scala 39:67]
          rdata <= _GEN_6;
        end else begin
          rdata <= _GEN_56;
        end
      end
    end
    if (io_cpu_req_valid) begin // @[Reg.scala 16:19]
      cpu_addr <= io_cpu_req_bits_addr; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[MMU.scala 75:22]
      state <= 4'h0; // @[MMU.scala 75:22]
    end else if (_T_27) begin // @[Conditional.scala 40:58]
      if (io_cpu_req_valid & _T_13 & MODE) begin // @[MMU.scala 116:62]
        state <= 4'h1; // @[MMU.scala 121:15]
      end
    end else if (_T_32) begin // @[Conditional.scala 39:67]
      state <= 4'h2; // @[MMU.scala 128:13]
    end else if (_T_33) begin // @[Conditional.scala 39:67]
      state <= _GEN_7;
    end else begin
      state <= _GEN_52;
    end
    if (reset) begin // @[MMU.scala 78:29]
      cacheReqAddr <= 32'h0; // @[MMU.scala 78:29]
    end else if (_T_27) begin // @[Conditional.scala 40:58]
      if (io_cpu_req_valid & _T_13 & MODE) begin // @[MMU.scala 116:62]
        cacheReqAddr <= io_cpu_req_bits_addr; // @[MMU.scala 118:22]
      end
    end
    if (reset) begin // @[MMU.scala 79:30]
      cacheReqData <= 32'h0; // @[MMU.scala 79:30]
    end else if (_T_27) begin // @[Conditional.scala 40:58]
      if (io_cpu_req_valid & _T_13 & MODE) begin // @[MMU.scala 116:62]
        cacheReqData <= io_cpu_req_bits_data; // @[MMU.scala 119:22]
      end
    end
    if (reset) begin // @[MMU.scala 80:30]
      cacheReqMask <= 4'h0; // @[MMU.scala 80:30]
    end else if (_T_27) begin // @[Conditional.scala 40:58]
      if (io_cpu_req_valid & _T_13 & MODE) begin // @[MMU.scala 116:62]
        cacheReqMask <= io_cpu_req_bits_mask; // @[MMU.scala 120:22]
      end
    end
    if (reset) begin // @[MMU.scala 97:26]
      pageFault <= 2'h0; // @[MMU.scala 97:26]
    end else if (_T_27) begin // @[Conditional.scala 40:58]
      if (clearPageFault_0) begin // @[MMU.scala 115:27]
        pageFault <= 2'h0; // @[MMU.scala 115:38]
      end
    end else if (!(_T_32)) begin // @[Conditional.scala 39:67]
      if (!(_T_33)) begin // @[Conditional.scala 39:67]
        pageFault <= _GEN_55;
      end
    end
    if (reset) begin // @[MMU.scala 108:28]
      cpuRespData <= 32'h0; // @[MMU.scala 108:28]
    end else if (!(_T_27)) begin // @[Conditional.scala 40:58]
      if (!(_T_32)) begin // @[Conditional.scala 39:67]
        if (!(_T_33)) begin // @[Conditional.scala 39:67]
          cpuRespData <= _GEN_59;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rdata = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cpu_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  cacheReqAddr = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  cacheReqData = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  cacheReqMask = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  pageFault = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  cpuRespData = _RAND_7[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RegMapper(
  input         clock,
  input         io_selector_req_valid,
  input  [31:0] io_selector_req_bits_addr,
  input  [31:0] io_selector_req_bits_data,
  input  [3:0]  io_selector_req_bits_mask,
  output        io_selector_resp_valid,
  output [31:0] io_selector_resp_bits_data,
  output        io_uart_req_valid,
  output [31:0] io_uart_req_bits_addr,
  output [31:0] io_uart_req_bits_data,
  input         io_uart_resp_valid,
  input  [31:0] io_uart_resp_bits_data,
  output        io_rtc_req_valid,
  output [31:0] io_rtc_req_bits_addr,
  output [31:0] io_rtc_req_bits_data,
  output [3:0]  io_rtc_req_bits_mask,
  input         io_rtc_resp_valid,
  input  [31:0] io_rtc_resp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] addr; // @[Reg.scala 15:16]
  wire [31:0] _T = io_selector_req_bits_addr & 32'hfffffff0; // @[RegMapper.scala 25:51]
  wire [31:0] _T_6 = addr & 32'hfffffff0; // @[RegMapper.scala 31:11]
  wire  _T_7 = 32'h10000000 == _T_6; // @[RegMapper.scala 31:11]
  wire  _T_9 = 32'h10010000 == _T_6; // @[RegMapper.scala 32:11]
  wire [31:0] _T_10 = _T_9 ? io_rtc_resp_bits_data : 32'h0; // @[Mux.scala 98:16]
  assign io_selector_resp_valid = _T_7 ? io_uart_resp_valid : _T_9 & io_rtc_resp_valid; // @[Mux.scala 98:16]
  assign io_selector_resp_bits_data = _T_7 ? io_uart_resp_bits_data : _T_10; // @[Mux.scala 98:16]
  assign io_uart_req_valid = 32'h10000000 == _T & io_selector_req_valid; // @[RegMapper.scala 25:71]
  assign io_uart_req_bits_addr = io_selector_req_bits_addr; // @[RegMapper.scala 24:20]
  assign io_uart_req_bits_data = io_selector_req_bits_data; // @[RegMapper.scala 24:20]
  assign io_rtc_req_valid = 32'h10010000 == _T & io_selector_req_valid; // @[RegMapper.scala 27:69]
  assign io_rtc_req_bits_addr = io_selector_req_bits_addr; // @[RegMapper.scala 26:19]
  assign io_rtc_req_bits_data = io_selector_req_bits_data; // @[RegMapper.scala 26:19]
  assign io_rtc_req_bits_mask = io_selector_req_bits_mask; // @[RegMapper.scala 26:19]
  always @(posedge clock) begin
    if (io_selector_req_valid) begin // @[Reg.scala 16:19]
      addr <= io_selector_req_bits_addr; // @[Reg.scala 16:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module DRAM(
  output        io_nasti_aw_ready,
  input         io_nasti_aw_valid,
  input  [31:0] io_nasti_aw_bits_addr,
  output        io_nasti_w_ready,
  input         io_nasti_w_valid,
  input  [31:0] io_nasti_w_bits_data,
  input         io_nasti_w_bits_last,
  input         io_nasti_b_ready,
  output        io_nasti_b_valid,
  output        io_nasti_ar_ready,
  input         io_nasti_ar_valid,
  input  [31:0] io_nasti_ar_bits_addr,
  input         io_nasti_r_ready,
  output        io_nasti_r_valid,
  output [31:0] io_nasti_r_bits_data,
  output        io_nasti_r_bits_last,
  output [31:0] io_AXI_s_axi_awaddr,
  output        io_AXI_s_axi_awvalid,
  input         io_AXI_s_axi_awready,
  output [31:0] io_AXI_s_axi_wdata,
  output        io_AXI_s_axi_wlast,
  output        io_AXI_s_axi_wvalid,
  input         io_AXI_s_axi_wready,
  input         io_AXI_s_axi_bvalid,
  output        io_AXI_s_axi_bready,
  output [31:0] io_AXI_s_axi_araddr,
  output        io_AXI_s_axi_arvalid,
  input         io_AXI_s_axi_arready,
  input  [31:0] io_AXI_s_axi_rdata,
  input         io_AXI_s_axi_rlast,
  input         io_AXI_s_axi_rvalid,
  output        io_AXI_s_axi_rready
);
  assign io_nasti_aw_ready = io_AXI_s_axi_awready; // @[DRAM.scala 54:21]
  assign io_nasti_w_ready = io_AXI_s_axi_wready; // @[DRAM.scala 59:20]
  assign io_nasti_b_valid = io_AXI_s_axi_bvalid; // @[DRAM.scala 62:20]
  assign io_nasti_ar_ready = io_AXI_s_axi_arready; // @[DRAM.scala 70:21]
  assign io_nasti_r_valid = io_AXI_s_axi_rvalid; // @[DRAM.scala 75:20]
  assign io_nasti_r_bits_data = io_AXI_s_axi_rdata; // @[DRAM.scala 72:24]
  assign io_nasti_r_bits_last = io_AXI_s_axi_rlast; // @[DRAM.scala 74:24]
  assign io_AXI_s_axi_awaddr = io_nasti_aw_bits_addr; // @[DRAM.scala 49:23]
  assign io_AXI_s_axi_awvalid = io_nasti_aw_valid; // @[DRAM.scala 53:24]
  assign io_AXI_s_axi_wdata = io_nasti_w_bits_data; // @[DRAM.scala 55:22]
  assign io_AXI_s_axi_wlast = io_nasti_w_bits_last; // @[DRAM.scala 57:22]
  assign io_AXI_s_axi_wvalid = io_nasti_w_valid; // @[DRAM.scala 58:23]
  assign io_AXI_s_axi_bready = io_nasti_b_ready; // @[DRAM.scala 63:23]
  assign io_AXI_s_axi_araddr = io_nasti_ar_bits_addr; // @[DRAM.scala 65:23]
  assign io_AXI_s_axi_arvalid = io_nasti_ar_valid; // @[DRAM.scala 69:24]
  assign io_AXI_s_axi_rready = io_nasti_r_ready; // @[DRAM.scala 76:23]
endmodule
module UartController(
  input         clock,
  input         reset,
  input         io__cpu_req_valid,
  input  [31:0] io__cpu_req_bits_addr,
  input  [31:0] io__cpu_req_bits_data,
  output        io__cpu_resp_valid,
  output [31:0] io__cpu_resp_bits_data,
  output        io__rxChannel_ready,
  input         io__rxChannel_valid,
  input  [7:0]  io__rxChannel_bits,
  input         io__txChannel_ready,
  output        io__txChannel_valid,
  output [7:0]  io__txChannel_bits,
  output        io_rxChannel_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Uart.scala 218:22]
  wire  is_READ_READ_STATE = state == 3'h1; // @[Uart.scala 220:34]
  wire  is_READ_WRITE_STATE = state == 3'h2; // @[Uart.scala 221:35]
  wire  is_READ_DATA = state == 3'h3; // @[Uart.scala 222:28]
  wire  _T_1 = is_READ_READ_STATE | is_READ_WRITE_STATE | is_READ_DATA; // @[Uart.scala 225:89]
  reg [31:0] rdata; // @[Reg.scala 15:16]
  reg [31:0] wdata; // @[Uart.scala 226:22]
  wire  _T_2 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire [2:0] _T_4 = 32'h10000000 == io__cpu_req_bits_addr ? 3'h1 : 3'h0; // @[Mux.scala 80:57]
  wire [2:0] _T_6 = 32'h10000004 == io__cpu_req_bits_addr ? 3'h3 : _T_4; // @[Mux.scala 80:57]
  wire [2:0] _T_8 = 32'h10000008 == io__cpu_req_bits_addr ? 3'h2 : _T_6; // @[Mux.scala 80:57]
  wire  _T_11 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_14 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_17 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_18 = io__rxChannel_ready & io__rxChannel_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_4 = _T_18 ? {{24'd0}, io__rxChannel_bits} : rdata; // @[Uart.scala 268:33 Uart.scala 269:31 Uart.scala 230:25]
  wire [2:0] _GEN_6 = _T_18 ? 3'h0 : state; // @[Uart.scala 268:33 Uart.scala 271:15 Uart.scala 218:22]
  wire  _T_19 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_21 = io__txChannel_ready & io__txChannel_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _GEN_7 = _T_21 ? 3'h0 : state; // @[Uart.scala 279:33 Uart.scala 280:15 Uart.scala 218:22]
  wire [7:0] _GEN_8 = _T_19 ? wdata[7:0] : 8'h0; // @[Conditional.scala 39:67 Uart.scala 277:25 Uart.scala 231:21]
  wire [2:0] _GEN_10 = _T_19 ? _GEN_7 : state; // @[Conditional.scala 39:67 Uart.scala 218:22]
  wire [31:0] _GEN_12 = _T_17 ? _GEN_4 : rdata; // @[Conditional.scala 39:67 Uart.scala 230:25]
  wire  _GEN_13 = _T_17 & _T_18; // @[Conditional.scala 39:67 Uart.scala 229:21]
  wire [2:0] _GEN_14 = _T_17 ? _GEN_6 : _GEN_10; // @[Conditional.scala 39:67]
  wire [7:0] _GEN_15 = _T_17 ? 8'h0 : _GEN_8; // @[Conditional.scala 39:67 Uart.scala 231:21]
  wire  _GEN_16 = _T_17 ? 1'h0 : _T_19; // @[Conditional.scala 39:67 Uart.scala 232:22]
  wire [31:0] _GEN_17 = _T_14 ? {{31'd0}, io__txChannel_ready} : _GEN_12; // @[Conditional.scala 39:67 Uart.scala 262:29]
  wire  _GEN_18 = _T_14 | _GEN_13; // @[Conditional.scala 39:67 Uart.scala 263:25]
  wire  _GEN_20 = _T_14 ? 1'h0 : _T_17; // @[Conditional.scala 39:67 Uart.scala 228:22]
  wire [7:0] _GEN_21 = _T_14 ? 8'h0 : _GEN_15; // @[Conditional.scala 39:67 Uart.scala 231:21]
  wire  _GEN_22 = _T_14 ? 1'h0 : _GEN_16; // @[Conditional.scala 39:67 Uart.scala 232:22]
  wire [31:0] _GEN_23 = _T_11 ? {{31'd0}, io__rxChannel_valid} : _GEN_17; // @[Conditional.scala 39:67 Uart.scala 256:29]
  wire  _GEN_24 = _T_11 | _GEN_18; // @[Conditional.scala 39:67 Uart.scala 257:25]
  wire  _GEN_26 = _T_11 ? 1'h0 : _GEN_20; // @[Conditional.scala 39:67 Uart.scala 228:22]
  wire [7:0] _GEN_27 = _T_11 ? 8'h0 : _GEN_21; // @[Conditional.scala 39:67 Uart.scala 231:21]
  wire  _GEN_28 = _T_11 ? 1'h0 : _GEN_22; // @[Conditional.scala 39:67 Uart.scala 232:22]
  assign io__cpu_resp_valid = _T_2 | _GEN_24; // @[Conditional.scala 40:58 Uart.scala 242:25]
  assign io__cpu_resp_bits_data = _T_2 ? rdata : _GEN_23; // @[Conditional.scala 40:58 Uart.scala 230:25]
  assign io__rxChannel_ready = _T_2 ? 1'h0 : _GEN_26; // @[Conditional.scala 40:58 Uart.scala 228:22]
  assign io__txChannel_valid = _T_2 ? 1'h0 : _GEN_28; // @[Conditional.scala 40:58 Uart.scala 232:22]
  assign io__txChannel_bits = _T_2 ? 8'h0 : _GEN_27; // @[Conditional.scala 40:58 Uart.scala 231:21]
  assign io_rxChannel_valid = io__rxChannel_valid;
  always @(posedge clock) begin
    if (reset) begin // @[Uart.scala 218:22]
      state <= 3'h0; // @[Uart.scala 218:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (io__cpu_req_valid) begin // @[Uart.scala 243:31]
        if (32'h1000000c == io__cpu_req_bits_addr) begin // @[Mux.scala 80:57]
          state <= 3'h4;
        end else begin
          state <= _T_8;
        end
      end
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      state <= 3'h0; // @[Uart.scala 258:13]
    end else if (_T_14) begin // @[Conditional.scala 39:67]
      state <= 3'h0; // @[Uart.scala 264:13]
    end else begin
      state <= _GEN_14;
    end
    if (_T_1) begin // @[Reg.scala 16:19]
      rdata <= io__cpu_resp_bits_data; // @[Reg.scala 16:23]
    end
    if (reset) begin // @[Uart.scala 226:22]
      wdata <= 32'h0; // @[Uart.scala 226:22]
    end else if (_T_2) begin // @[Conditional.scala 40:58]
      if (io__cpu_req_valid) begin // @[Uart.scala 243:31]
        wdata <= io__cpu_req_bits_data; // @[Uart.scala 245:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  rdata = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  wdata = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Tx(
  input        clock,
  input        reset,
  output       io_txd,
  output       io_channel_ready,
  input        io_channel_valid,
  input  [7:0] io_channel_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  state; // @[Uart.scala 32:22]
  reg [10:0] shiftReg; // @[Uart.scala 36:25]
  reg [7:0] baud_count; // @[Counter.scala 60:40]
  wire  wrap_wrap = baud_count == 8'hc1; // @[Counter.scala 72:24]
  wire [7:0] _wrap_value_T_1 = baud_count + 8'h1; // @[Counter.scala 76:24]
  wire  baud_wrap_out = state & wrap_wrap; // @[Counter.scala 118:17 Counter.scala 118:24]
  reg [3:0] bit_count; // @[Counter.scala 60:40]
  wire  wrap_wrap_1 = bit_count == 4'ha; // @[Counter.scala 72:24]
  wire [3:0] _wrap_value_T_3 = bit_count + 4'h1; // @[Counter.scala 76:24]
  wire  bit_wrap_out = baud_wrap_out & wrap_wrap_1; // @[Counter.scala 118:17 Counter.scala 118:24]
  wire  _T_1 = ~state; // @[Uart.scala 43:29]
  wire  _T_3 = io_channel_ready & io_channel_valid; // @[Decoupled.scala 40:37]
  wire [10:0] _T_4 = {2'h3,io_channel_bits,1'h0}; // @[Cat.scala 30:58]
  wire [10:0] _GEN_6 = _T_3 ? _T_4 : shiftReg; // @[Uart.scala 47:27 Uart.scala 48:14 Uart.scala 36:25]
  wire [9:0] lo = shiftReg[10:1]; // @[Uart.scala 52:28]
  wire [10:0] _T_7 = {1'h1,lo}; // @[Cat.scala 30:58]
  wire  _GEN_9 = _T_3 | state; // @[Uart.scala 60:31 Uart.scala 61:15 Uart.scala 32:22]
  assign io_txd = shiftReg[0]; // @[Uart.scala 44:21]
  assign io_channel_ready = ~state; // @[Uart.scala 43:29]
  always @(posedge clock) begin
    if (reset) begin // @[Uart.scala 32:22]
      state <= 1'h0; // @[Uart.scala 32:22]
    end else if (_T_1) begin // @[Conditional.scala 40:58]
      state <= _GEN_9;
    end else if (state) begin // @[Conditional.scala 39:67]
      if (bit_wrap_out) begin // @[Uart.scala 65:26]
        state <= 1'h0; // @[Uart.scala 66:15]
      end
    end
    if (reset) begin // @[Uart.scala 36:25]
      shiftReg <= 11'h7ff; // @[Uart.scala 36:25]
    end else if (state) begin // @[Uart.scala 50:26]
      if (baud_wrap_out) begin // @[Uart.scala 51:25]
        shiftReg <= _T_7; // @[Uart.scala 53:16]
      end else begin
        shiftReg <= _GEN_6;
      end
    end else begin
      shiftReg <= _GEN_6;
    end
    if (reset) begin // @[Counter.scala 60:40]
      baud_count <= 8'h0; // @[Counter.scala 60:40]
    end else if (state) begin // @[Counter.scala 118:17]
      if (wrap_wrap) begin // @[Counter.scala 86:20]
        baud_count <= 8'h0; // @[Counter.scala 86:28]
      end else begin
        baud_count <= _wrap_value_T_1; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      bit_count <= 4'h0; // @[Counter.scala 60:40]
    end else if (baud_wrap_out) begin // @[Counter.scala 118:17]
      if (wrap_wrap_1) begin // @[Counter.scala 86:20]
        bit_count <= 4'h0; // @[Counter.scala 86:28]
      end else begin
        bit_count <= _wrap_value_T_3; // @[Counter.scala 76:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  shiftReg = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  baud_count = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  bit_count = _RAND_3[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Buffer(
  input        clock,
  input        reset,
  output       io_in_ready,
  input        io_in_valid,
  input  [7:0] io_in_bits,
  input        io_out_ready,
  output       io_out_valid,
  output [7:0] io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  state; // @[Uart.scala 79:22]
  reg [7:0] data; // @[Uart.scala 80:21]
  wire  _T = ~state; // @[Uart.scala 82:24]
  wire  _T_3 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_1 = _T_3 | state; // @[Uart.scala 88:26 Uart.scala 90:15 Uart.scala 79:22]
  wire  _T_5 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = ~state; // @[Uart.scala 82:24]
  assign io_out_valid = state; // @[Uart.scala 83:25]
  assign io_out_bits = data; // @[Uart.scala 84:15]
  always @(posedge clock) begin
    if (reset) begin // @[Uart.scala 79:22]
      state <= 1'h0; // @[Uart.scala 79:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      state <= _GEN_1;
    end else if (state) begin // @[Conditional.scala 39:67]
      if (_T_5) begin // @[Uart.scala 94:27]
        state <= 1'h0; // @[Uart.scala 95:15]
      end
    end
    if (reset) begin // @[Uart.scala 80:21]
      data <= 8'h0; // @[Uart.scala 80:21]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (_T_3) begin // @[Uart.scala 88:26]
        data <= io_in_bits; // @[Uart.scala 89:14]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  data = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BufferedTx(
  input        clock,
  input        reset,
  output       io_txd,
  output       io_channel_ready,
  input        io_channel_valid,
  input  [7:0] io_channel_bits
);
  wire  tx_clock; // @[Uart.scala 135:18]
  wire  tx_reset; // @[Uart.scala 135:18]
  wire  tx_io_txd; // @[Uart.scala 135:18]
  wire  tx_io_channel_ready; // @[Uart.scala 135:18]
  wire  tx_io_channel_valid; // @[Uart.scala 135:18]
  wire [7:0] tx_io_channel_bits; // @[Uart.scala 135:18]
  wire  buf__clock; // @[Uart.scala 136:19]
  wire  buf__reset; // @[Uart.scala 136:19]
  wire  buf__io_in_ready; // @[Uart.scala 136:19]
  wire  buf__io_in_valid; // @[Uart.scala 136:19]
  wire [7:0] buf__io_in_bits; // @[Uart.scala 136:19]
  wire  buf__io_out_ready; // @[Uart.scala 136:19]
  wire  buf__io_out_valid; // @[Uart.scala 136:19]
  wire [7:0] buf__io_out_bits; // @[Uart.scala 136:19]
  Tx tx ( // @[Uart.scala 135:18]
    .clock(tx_clock),
    .reset(tx_reset),
    .io_txd(tx_io_txd),
    .io_channel_ready(tx_io_channel_ready),
    .io_channel_valid(tx_io_channel_valid),
    .io_channel_bits(tx_io_channel_bits)
  );
  Buffer buf_ ( // @[Uart.scala 136:19]
    .clock(buf__clock),
    .reset(buf__reset),
    .io_in_ready(buf__io_in_ready),
    .io_in_valid(buf__io_in_valid),
    .io_in_bits(buf__io_in_bits),
    .io_out_ready(buf__io_out_ready),
    .io_out_valid(buf__io_out_valid),
    .io_out_bits(buf__io_out_bits)
  );
  assign io_txd = tx_io_txd; // @[Uart.scala 140:10]
  assign io_channel_ready = buf__io_in_ready; // @[Uart.scala 138:13]
  assign tx_clock = clock;
  assign tx_reset = reset;
  assign tx_io_channel_valid = buf__io_out_valid; // @[Uart.scala 139:17]
  assign tx_io_channel_bits = buf__io_out_bits; // @[Uart.scala 139:17]
  assign buf__clock = clock;
  assign buf__reset = reset;
  assign buf__io_in_valid = io_channel_valid; // @[Uart.scala 138:13]
  assign buf__io_in_bits = io_channel_bits; // @[Uart.scala 138:13]
  assign buf__io_out_ready = tx_io_channel_ready; // @[Uart.scala 139:17]
endmodule
module Rx(
  input        clock,
  input        reset,
  input        io_rxd,
  output       io_channel_valid,
  output [7:0] io_channel_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] shiftReg; // @[Uart.scala 149:25]
  reg [1:0] state; // @[Uart.scala 151:22]
  wire  _T = state == 2'h1; // @[Uart.scala 157:53]
  reg [8:0] first_count; // @[Counter.scala 60:40]
  wire  wrap_wrap = first_count == 9'h122; // @[Counter.scala 72:24]
  wire [8:0] _wrap_value_T_1 = first_count + 9'h1; // @[Counter.scala 76:24]
  wire  first_wrap_out = _T & wrap_wrap; // @[Counter.scala 118:17 Counter.scala 118:24]
  wire  _T_3 = state == 2'h2 | state == 2'h3; // @[Uart.scala 158:65]
  reg [7:0] baud_count; // @[Counter.scala 60:40]
  wire  wrap_wrap_1 = baud_count == 8'hc1; // @[Counter.scala 72:24]
  wire [7:0] _wrap_value_T_3 = baud_count + 8'h1; // @[Counter.scala 76:24]
  wire  baud_wrap_out = _T_3 & wrap_wrap_1; // @[Counter.scala 118:17 Counter.scala 118:24]
  wire  _T_4 = baud_wrap_out | first_wrap_out; // @[Uart.scala 159:58]
  wire  _T_6 = (baud_wrap_out | first_wrap_out) & state != 2'h3; // @[Uart.scala 159:77]
  reg [2:0] bit_count; // @[Counter.scala 60:40]
  wire  wrap_wrap_2 = bit_count == 3'h7; // @[Counter.scala 72:24]
  wire [2:0] _wrap_value_T_5 = bit_count + 3'h1; // @[Counter.scala 76:24]
  wire  bit_wrap_out = _T_6 & wrap_wrap_2; // @[Counter.scala 118:17 Counter.scala 118:24]
  wire [6:0] lo = shiftReg[7:1]; // @[Uart.scala 163:38]
  wire [7:0] _T_8 = {io_rxd,lo}; // @[Cat.scala 30:58]
  reg  REG; // @[Uart.scala 168:30]
  wire  _T_9 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_11 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_12 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_11 = bit_wrap_out ? 2'h3 : state; // @[Uart.scala 183:26 Uart.scala 184:15 Uart.scala 151:22]
  wire  _T_13 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_12 = baud_wrap_out ? 2'h0 : state; // @[Uart.scala 188:27 Uart.scala 189:15 Uart.scala 151:22]
  wire [1:0] _GEN_13 = _T_13 ? _GEN_12 : state; // @[Conditional.scala 39:67 Uart.scala 151:22]
  assign io_channel_valid = REG; // @[Uart.scala 168:20]
  assign io_channel_bits = shiftReg; // @[Uart.scala 167:19]
  always @(posedge clock) begin
    if (reset) begin // @[Uart.scala 149:25]
      shiftReg <= 8'h0; // @[Uart.scala 149:25]
    end else if (_T_4) begin // @[Uart.scala 162:41]
      shiftReg <= _T_8; // @[Uart.scala 163:14]
    end
    if (reset) begin // @[Uart.scala 151:22]
      state <= 2'h0; // @[Uart.scala 151:22]
    end else if (_T_9) begin // @[Conditional.scala 40:58]
      if (~io_rxd) begin // @[Uart.scala 173:28]
        state <= 2'h1; // @[Uart.scala 174:15]
      end
    end else if (_T_11) begin // @[Conditional.scala 39:67]
      if (first_wrap_out) begin // @[Uart.scala 178:28]
        state <= 2'h2; // @[Uart.scala 179:15]
      end
    end else if (_T_12) begin // @[Conditional.scala 39:67]
      state <= _GEN_11;
    end else begin
      state <= _GEN_13;
    end
    if (reset) begin // @[Counter.scala 60:40]
      first_count <= 9'h0; // @[Counter.scala 60:40]
    end else if (_T) begin // @[Counter.scala 118:17]
      if (wrap_wrap) begin // @[Counter.scala 86:20]
        first_count <= 9'h0; // @[Counter.scala 86:28]
      end else begin
        first_count <= _wrap_value_T_1; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      baud_count <= 8'h0; // @[Counter.scala 60:40]
    end else if (_T_3) begin // @[Counter.scala 118:17]
      if (wrap_wrap_1) begin // @[Counter.scala 86:20]
        baud_count <= 8'h0; // @[Counter.scala 86:28]
      end else begin
        baud_count <= _wrap_value_T_3; // @[Counter.scala 76:15]
      end
    end
    if (reset) begin // @[Counter.scala 60:40]
      bit_count <= 3'h0; // @[Counter.scala 60:40]
    end else if (_T_6) begin // @[Counter.scala 118:17]
      bit_count <= _wrap_value_T_5; // @[Counter.scala 76:15]
    end
    REG <= _T_6 & wrap_wrap_2; // @[Counter.scala 118:17 Counter.scala 118:24]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  shiftReg = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  first_count = _RAND_2[8:0];
  _RAND_3 = {1{`RANDOM}};
  baud_count = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  bit_count = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  REG = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BufferedRx(
  input        clock,
  input        reset,
  input        io_rxd,
  input        io_channel_ready,
  output       io_channel_valid,
  output [7:0] io_channel_bits
);
  wire  rx_clock; // @[Uart.scala 201:18]
  wire  rx_reset; // @[Uart.scala 201:18]
  wire  rx_io_rxd; // @[Uart.scala 201:18]
  wire  rx_io_channel_valid; // @[Uart.scala 201:18]
  wire [7:0] rx_io_channel_bits; // @[Uart.scala 201:18]
  wire  buf__clock; // @[Uart.scala 202:19]
  wire  buf__reset; // @[Uart.scala 202:19]
  wire  buf__io_in_ready; // @[Uart.scala 202:19]
  wire  buf__io_in_valid; // @[Uart.scala 202:19]
  wire [7:0] buf__io_in_bits; // @[Uart.scala 202:19]
  wire  buf__io_out_ready; // @[Uart.scala 202:19]
  wire  buf__io_out_valid; // @[Uart.scala 202:19]
  wire [7:0] buf__io_out_bits; // @[Uart.scala 202:19]
  Rx rx ( // @[Uart.scala 201:18]
    .clock(rx_clock),
    .reset(rx_reset),
    .io_rxd(rx_io_rxd),
    .io_channel_valid(rx_io_channel_valid),
    .io_channel_bits(rx_io_channel_bits)
  );
  Buffer buf_ ( // @[Uart.scala 202:19]
    .clock(buf__clock),
    .reset(buf__reset),
    .io_in_ready(buf__io_in_ready),
    .io_in_valid(buf__io_in_valid),
    .io_in_bits(buf__io_in_bits),
    .io_out_ready(buf__io_out_ready),
    .io_out_valid(buf__io_out_valid),
    .io_out_bits(buf__io_out_bits)
  );
  assign io_channel_valid = buf__io_out_valid; // @[Uart.scala 206:14]
  assign io_channel_bits = buf__io_out_bits; // @[Uart.scala 206:14]
  assign rx_clock = clock;
  assign rx_reset = reset;
  assign rx_io_rxd = io_rxd; // @[Uart.scala 204:10]
  assign buf__clock = clock;
  assign buf__reset = reset;
  assign buf__io_in_valid = rx_io_channel_valid; // @[Uart.scala 205:13]
  assign buf__io_in_bits = rx_io_channel_bits; // @[Uart.scala 205:13]
  assign buf__io_out_ready = io_channel_ready; // @[Uart.scala 206:14]
endmodule
module Uart(
  input        clock,
  input        reset,
  input        io_rxd,
  output       io_txd,
  input        io_rxChannel_ready,
  output       io_rxChannel_valid,
  output [7:0] io_rxChannel_bits,
  output       io_txChannel_ready,
  input        io_txChannel_valid,
  input  [7:0] io_txChannel_bits
);
  wire  tx_clock; // @[Uart.scala 294:18]
  wire  tx_reset; // @[Uart.scala 294:18]
  wire  tx_io_txd; // @[Uart.scala 294:18]
  wire  tx_io_channel_ready; // @[Uart.scala 294:18]
  wire  tx_io_channel_valid; // @[Uart.scala 294:18]
  wire [7:0] tx_io_channel_bits; // @[Uart.scala 294:18]
  wire  rx_clock; // @[Uart.scala 295:18]
  wire  rx_reset; // @[Uart.scala 295:18]
  wire  rx_io_rxd; // @[Uart.scala 295:18]
  wire  rx_io_channel_ready; // @[Uart.scala 295:18]
  wire  rx_io_channel_valid; // @[Uart.scala 295:18]
  wire [7:0] rx_io_channel_bits; // @[Uart.scala 295:18]
  BufferedTx tx ( // @[Uart.scala 294:18]
    .clock(tx_clock),
    .reset(tx_reset),
    .io_txd(tx_io_txd),
    .io_channel_ready(tx_io_channel_ready),
    .io_channel_valid(tx_io_channel_valid),
    .io_channel_bits(tx_io_channel_bits)
  );
  BufferedRx rx ( // @[Uart.scala 295:18]
    .clock(rx_clock),
    .reset(rx_reset),
    .io_rxd(rx_io_rxd),
    .io_channel_ready(rx_io_channel_ready),
    .io_channel_valid(rx_io_channel_valid),
    .io_channel_bits(rx_io_channel_bits)
  );
  assign io_txd = tx_io_txd; // @[Uart.scala 299:13]
  assign io_rxChannel_valid = rx_io_channel_valid; // @[Uart.scala 298:17]
  assign io_rxChannel_bits = rx_io_channel_bits; // @[Uart.scala 298:17]
  assign io_txChannel_ready = tx_io_channel_ready; // @[Uart.scala 297:17]
  assign tx_clock = clock;
  assign tx_reset = reset;
  assign tx_io_channel_valid = io_txChannel_valid; // @[Uart.scala 297:17]
  assign tx_io_channel_bits = io_txChannel_bits; // @[Uart.scala 297:17]
  assign rx_clock = clock;
  assign rx_reset = reset;
  assign rx_io_rxd = io_rxd; // @[Uart.scala 300:13]
  assign rx_io_channel_ready = io_rxChannel_ready; // @[Uart.scala 298:17]
endmodule
module RTC(
  input         clock,
  input         reset,
  input         io_req_valid,
  input  [31:0] io_req_bits_addr,
  input  [31:0] io_req_bits_data,
  input  [3:0]  io_req_bits_mask,
  output        io_resp_valid,
  output [31:0] io_resp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] time_; // @[RTC.scala 17:21]
  reg [31:0] timeh; // @[RTC.scala 18:22]
  reg [1:0] state; // @[RTC.scala 19:22]
  reg [3:0] mask; // @[RTC.scala 21:21]
  reg [31:0] data; // @[RTC.scala 22:21]
  reg [31:0] cntReg; // @[RTC.scala 29:23]
  wire [31:0] _T_1 = cntReg + 32'h1; // @[RTC.scala 31:20]
  wire [31:0] _T_4 = time_ + 32'h1; // @[RTC.scala 34:18]
  wire [31:0] _T_7 = timeh + 32'h1; // @[RTC.scala 36:38]
  wire [31:0] _GEN_0 = &time_ ? _T_7 : timeh; // @[RTC.scala 36:21 RTC.scala 36:29 RTC.scala 18:22]
  wire [31:0] _GEN_2 = cntReg == 32'h98967f ? _T_4 : time_; // @[RTC.scala 32:27 RTC.scala 34:10 RTC.scala 17:21]
  wire [31:0] _GEN_3 = cntReg == 32'h98967f ? _GEN_0 : timeh; // @[RTC.scala 32:27 RTC.scala 18:22]
  wire  _T_8 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire [31:0] _T_9 = io_req_bits_addr & 32'h1fffffff; // @[RTC.scala 48:29]
  wire  _T_10 = 32'h10001000 == _T_9; // @[RTC.scala 48:29]
  wire  _T_12 = 32'h10001004 == _T_9; // @[RTC.scala 49:29]
  wire [1:0] _T_13 = _T_12 ? 2'h2 : 2'h0; // @[Mux.scala 98:16]
  wire  _T_15 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_17 = ~(|mask); // @[RTC.scala 54:14]
  wire [31:0] _GEN_8 = ~(|mask) ? time_ : 32'h0; // @[RTC.scala 54:26 RTC.scala 55:30 RTC.scala 24:21]
  wire  _T_18 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_11 = _T_17 ? timeh : 32'h0; // @[RTC.scala 63:24 RTC.scala 64:27 RTC.scala 24:21]
  wire [31:0] _GEN_13 = _T_17 ? _GEN_3 : data; // @[RTC.scala 63:24 RTC.scala 67:15]
  wire [31:0] _GEN_14 = _T_18 ? _GEN_11 : 32'h0; // @[Conditional.scala 39:67 RTC.scala 24:21]
  wire  _GEN_15 = _T_18 & _T_17; // @[Conditional.scala 39:67 RTC.scala 25:17]
  wire [31:0] _GEN_18 = _T_15 ? _GEN_8 : _GEN_14; // @[Conditional.scala 39:67]
  wire  _GEN_19 = _T_15 ? _T_17 : _GEN_15; // @[Conditional.scala 39:67]
  assign io_resp_valid = _T_8 | _GEN_19; // @[Conditional.scala 40:58 RTC.scala 42:21]
  assign io_resp_bits_data = _T_8 ? 32'h0 : _GEN_18; // @[Conditional.scala 40:58 RTC.scala 24:21]
  always @(posedge clock) begin
    if (reset) begin // @[RTC.scala 17:21]
      time_ <= 32'h0; // @[RTC.scala 17:21]
    end else if (_T_8) begin // @[Conditional.scala 40:58]
      time_ <= _GEN_2;
    end else if (_T_15) begin // @[Conditional.scala 39:67]
      if (~(|mask)) begin // @[RTC.scala 54:26]
        time_ <= _GEN_2;
      end else begin
        time_ <= data; // @[RTC.scala 58:16]
      end
    end else begin
      time_ <= _GEN_2;
    end
    if (reset) begin // @[RTC.scala 18:22]
      timeh <= 32'h0; // @[RTC.scala 18:22]
    end else if (_T_8) begin // @[Conditional.scala 40:58]
      timeh <= _GEN_3;
    end else if (_T_15) begin // @[Conditional.scala 39:67]
      timeh <= _GEN_3;
    end else if (_T_18) begin // @[Conditional.scala 39:67]
      timeh <= _GEN_13;
    end else begin
      timeh <= _GEN_3;
    end
    if (reset) begin // @[RTC.scala 19:22]
      state <= 2'h0; // @[RTC.scala 19:22]
    end else if (_T_8) begin // @[Conditional.scala 40:58]
      if (io_req_valid) begin // @[RTC.scala 43:26]
        if (_T_10) begin // @[Mux.scala 98:16]
          state <= 2'h1;
        end else begin
          state <= _T_13;
        end
      end
    end else if (_T_15) begin // @[Conditional.scala 39:67]
      state <= 2'h0; // @[RTC.scala 60:13]
    end else if (_T_18) begin // @[Conditional.scala 39:67]
      state <= 2'h0; // @[RTC.scala 69:13]
    end
    if (reset) begin // @[RTC.scala 21:21]
      mask <= 4'h0; // @[RTC.scala 21:21]
    end else if (_T_8) begin // @[Conditional.scala 40:58]
      if (io_req_valid) begin // @[RTC.scala 43:26]
        mask <= io_req_bits_mask; // @[RTC.scala 45:14]
      end
    end
    if (reset) begin // @[RTC.scala 22:21]
      data <= 32'h0; // @[RTC.scala 22:21]
    end else if (_T_8) begin // @[Conditional.scala 40:58]
      if (io_req_valid) begin // @[RTC.scala 43:26]
        data <= io_req_bits_data; // @[RTC.scala 46:14]
      end
    end
    if (reset) begin // @[RTC.scala 29:23]
      cntReg <= 32'h0; // @[RTC.scala 29:23]
    end else if (cntReg == 32'h98967f) begin // @[RTC.scala 32:27]
      cntReg <= 32'h0; // @[RTC.scala 33:12]
    end else begin
      cntReg <= _T_1; // @[RTC.scala 31:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  time_ = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  timeh = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  mask = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  data = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  cntReg = _RAND_5[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Tile(
  input         clock,
  input         reset,
  output [3:0]  io_AXI_s_axi_awid,
  output [31:0] io_AXI_s_axi_awaddr,
  output [7:0]  io_AXI_s_axi_awlen,
  output [2:0]  io_AXI_s_axi_awsize,
  output [1:0]  io_AXI_s_axi_awburst,
  output        io_AXI_s_axi_awvalid,
  input         io_AXI_s_axi_awready,
  output [31:0] io_AXI_s_axi_wdata,
  output [7:0]  io_AXI_s_axi_wstrb,
  output        io_AXI_s_axi_wlast,
  output        io_AXI_s_axi_wvalid,
  input         io_AXI_s_axi_wready,
  input  [3:0]  io_AXI_s_axi_bid,
  input  [1:0]  io_AXI_s_axi_bresp,
  input         io_AXI_s_axi_bvalid,
  output        io_AXI_s_axi_bready,
  output [3:0]  io_AXI_s_axi_arid,
  output [31:0] io_AXI_s_axi_araddr,
  output [7:0]  io_AXI_s_axi_arlen,
  output [2:0]  io_AXI_s_axi_arsize,
  output [1:0]  io_AXI_s_axi_arburst,
  output        io_AXI_s_axi_arvalid,
  input         io_AXI_s_axi_arready,
  input  [3:0]  io_AXI_s_axi_rid,
  input  [31:0] io_AXI_s_axi_rdata,
  input  [1:0]  io_AXI_s_axi_rresp,
  input         io_AXI_s_axi_rlast,
  input         io_AXI_s_axi_rvalid,
  output        io_AXI_s_axi_rready,
  output        io_txd,
  input         io_rxd
);
  wire  dfc_table_clock; // @[Tile.scala 120:25]
  wire  dfc_table_reset; // @[Tile.scala 120:25]
  wire  dfc_table_io_cpu1_w_data_valid; // @[Tile.scala 120:25]
  wire [31:0] dfc_table_io_cpu1_w_data_bits_listenAddr; // @[Tile.scala 120:25]
  wire [15:0] dfc_table_io_cpu1_w_data_bits_wPid; // @[Tile.scala 120:25]
  wire  dfc_table_io_cpu1_l_data_valid; // @[Tile.scala 120:25]
  wire [31:0] dfc_table_io_cpu1_l_data_bits_listenAddr; // @[Tile.scala 120:25]
  wire  dfc_table_io_cpu1_e_data_ready; // @[Tile.scala 120:25]
  wire  dfc_table_io_cpu1_e_data_valid; // @[Tile.scala 120:25]
  wire [15:0] dfc_table_io_cpu1_e_data_bits_pid; // @[Tile.scala 120:25]
  wire  dfc_table_io_cpu_f_data_valid; // @[Tile.scala 120:25]
  wire  dfc_table_io_cpu_f_data_bits_full_sig; // @[Tile.scala 120:25]
  wire  core_clock; // @[Tile.scala 125:20]
  wire  core_reset; // @[Tile.scala 125:20]
  wire  core_io_icache_req_valid; // @[Tile.scala 125:20]
  wire [31:0] core_io_icache_req_bits_addr; // @[Tile.scala 125:20]
  wire  core_io_icache_resp_valid; // @[Tile.scala 125:20]
  wire [31:0] core_io_icache_resp_bits_data; // @[Tile.scala 125:20]
  wire  core_io_dcache_abort; // @[Tile.scala 125:20]
  wire  core_io_dcache_req_valid; // @[Tile.scala 125:20]
  wire [31:0] core_io_dcache_req_bits_addr; // @[Tile.scala 125:20]
  wire [31:0] core_io_dcache_req_bits_data; // @[Tile.scala 125:20]
  wire [3:0] core_io_dcache_req_bits_mask; // @[Tile.scala 125:20]
  wire  core_io_dcache_resp_valid; // @[Tile.scala 125:20]
  wire [31:0] core_io_dcache_resp_bits_data; // @[Tile.scala 125:20]
  wire  core_io_table_w_data_valid; // @[Tile.scala 125:20]
  wire [31:0] core_io_table_w_data_bits_listenAddr; // @[Tile.scala 125:20]
  wire [15:0] core_io_table_w_data_bits_wPid; // @[Tile.scala 125:20]
  wire  core_io_table_l_data_valid; // @[Tile.scala 125:20]
  wire [31:0] core_io_table_l_data_bits_listenAddr; // @[Tile.scala 125:20]
  wire  core_io_table_e_data_ready; // @[Tile.scala 125:20]
  wire  core_io_table_e_data_valid; // @[Tile.scala 125:20]
  wire [15:0] core_io_table_e_data_bits_pid; // @[Tile.scala 125:20]
  wire  core_io_table_f_data_valid; // @[Tile.scala 125:20]
  wire  core_io_table_f_data_bits_full_sig; // @[Tile.scala 125:20]
  wire  core_io_rxChannel_valid; // @[Tile.scala 125:20]
  wire [1:0] core_pageFault; // @[Tile.scala 125:20]
  wire  core_io_vmSwitch; // @[Tile.scala 125:20]
  wire [31:0] core_io_in; // @[Tile.scala 125:20]
  wire  core_clearPageFault; // @[Tile.scala 125:20]
  wire [1:0] core_pageFault_0; // @[Tile.scala 125:20]
  wire [31:0] core_satp; // @[Tile.scala 125:20]
  wire  icache_clock; // @[Tile.scala 126:22]
  wire  icache_reset; // @[Tile.scala 126:22]
  wire  icache_io_cpu_abort; // @[Tile.scala 126:22]
  wire  icache_io_cpu_req_valid; // @[Tile.scala 126:22]
  wire [31:0] icache_io_cpu_req_bits_addr; // @[Tile.scala 126:22]
  wire [31:0] icache_io_cpu_req_bits_data; // @[Tile.scala 126:22]
  wire [3:0] icache_io_cpu_req_bits_mask; // @[Tile.scala 126:22]
  wire  icache_io_cpu_resp_valid; // @[Tile.scala 126:22]
  wire [31:0] icache_io_cpu_resp_bits_data; // @[Tile.scala 126:22]
  wire  icache_io_nasti_aw_ready; // @[Tile.scala 126:22]
  wire  icache_io_nasti_aw_valid; // @[Tile.scala 126:22]
  wire [31:0] icache_io_nasti_aw_bits_addr; // @[Tile.scala 126:22]
  wire  icache_io_nasti_w_ready; // @[Tile.scala 126:22]
  wire  icache_io_nasti_w_valid; // @[Tile.scala 126:22]
  wire [31:0] icache_io_nasti_w_bits_data; // @[Tile.scala 126:22]
  wire  icache_io_nasti_w_bits_last; // @[Tile.scala 126:22]
  wire  icache_io_nasti_b_ready; // @[Tile.scala 126:22]
  wire  icache_io_nasti_b_valid; // @[Tile.scala 126:22]
  wire  icache_io_nasti_ar_ready; // @[Tile.scala 126:22]
  wire  icache_io_nasti_ar_valid; // @[Tile.scala 126:22]
  wire [31:0] icache_io_nasti_ar_bits_addr; // @[Tile.scala 126:22]
  wire  icache_io_nasti_r_ready; // @[Tile.scala 126:22]
  wire  icache_io_nasti_r_valid; // @[Tile.scala 126:22]
  wire [31:0] icache_io_nasti_r_bits_data; // @[Tile.scala 126:22]
  wire  dcache_clock; // @[Tile.scala 127:22]
  wire  dcache_reset; // @[Tile.scala 127:22]
  wire  dcache_io_cpu_abort; // @[Tile.scala 127:22]
  wire  dcache_io_cpu_req_valid; // @[Tile.scala 127:22]
  wire [31:0] dcache_io_cpu_req_bits_addr; // @[Tile.scala 127:22]
  wire [31:0] dcache_io_cpu_req_bits_data; // @[Tile.scala 127:22]
  wire [3:0] dcache_io_cpu_req_bits_mask; // @[Tile.scala 127:22]
  wire  dcache_io_cpu_resp_valid; // @[Tile.scala 127:22]
  wire [31:0] dcache_io_cpu_resp_bits_data; // @[Tile.scala 127:22]
  wire  dcache_io_nasti_aw_ready; // @[Tile.scala 127:22]
  wire  dcache_io_nasti_aw_valid; // @[Tile.scala 127:22]
  wire [31:0] dcache_io_nasti_aw_bits_addr; // @[Tile.scala 127:22]
  wire  dcache_io_nasti_w_ready; // @[Tile.scala 127:22]
  wire  dcache_io_nasti_w_valid; // @[Tile.scala 127:22]
  wire [31:0] dcache_io_nasti_w_bits_data; // @[Tile.scala 127:22]
  wire  dcache_io_nasti_w_bits_last; // @[Tile.scala 127:22]
  wire  dcache_io_nasti_b_ready; // @[Tile.scala 127:22]
  wire  dcache_io_nasti_b_valid; // @[Tile.scala 127:22]
  wire  dcache_io_nasti_ar_ready; // @[Tile.scala 127:22]
  wire  dcache_io_nasti_ar_valid; // @[Tile.scala 127:22]
  wire [31:0] dcache_io_nasti_ar_bits_addr; // @[Tile.scala 127:22]
  wire  dcache_io_nasti_r_ready; // @[Tile.scala 127:22]
  wire  dcache_io_nasti_r_valid; // @[Tile.scala 127:22]
  wire [31:0] dcache_io_nasti_r_bits_data; // @[Tile.scala 127:22]
  wire  arb_clock; // @[Tile.scala 128:19]
  wire  arb_reset; // @[Tile.scala 128:19]
  wire  arb_io_icache_ar_ready; // @[Tile.scala 128:19]
  wire  arb_io_icache_ar_valid; // @[Tile.scala 128:19]
  wire [31:0] arb_io_icache_ar_bits_addr; // @[Tile.scala 128:19]
  wire  arb_io_icache_r_ready; // @[Tile.scala 128:19]
  wire  arb_io_icache_r_valid; // @[Tile.scala 128:19]
  wire [31:0] arb_io_icache_r_bits_data; // @[Tile.scala 128:19]
  wire  arb_io_dcache_aw_ready; // @[Tile.scala 128:19]
  wire  arb_io_dcache_aw_valid; // @[Tile.scala 128:19]
  wire [31:0] arb_io_dcache_aw_bits_addr; // @[Tile.scala 128:19]
  wire  arb_io_dcache_w_ready; // @[Tile.scala 128:19]
  wire  arb_io_dcache_w_valid; // @[Tile.scala 128:19]
  wire [31:0] arb_io_dcache_w_bits_data; // @[Tile.scala 128:19]
  wire  arb_io_dcache_w_bits_last; // @[Tile.scala 128:19]
  wire  arb_io_dcache_b_ready; // @[Tile.scala 128:19]
  wire  arb_io_dcache_b_valid; // @[Tile.scala 128:19]
  wire  arb_io_dcache_ar_ready; // @[Tile.scala 128:19]
  wire  arb_io_dcache_ar_valid; // @[Tile.scala 128:19]
  wire [31:0] arb_io_dcache_ar_bits_addr; // @[Tile.scala 128:19]
  wire  arb_io_dcache_r_ready; // @[Tile.scala 128:19]
  wire  arb_io_dcache_r_valid; // @[Tile.scala 128:19]
  wire [31:0] arb_io_dcache_r_bits_data; // @[Tile.scala 128:19]
  wire  arb_io_nasti_aw_ready; // @[Tile.scala 128:19]
  wire  arb_io_nasti_aw_valid; // @[Tile.scala 128:19]
  wire [31:0] arb_io_nasti_aw_bits_addr; // @[Tile.scala 128:19]
  wire  arb_io_nasti_w_ready; // @[Tile.scala 128:19]
  wire  arb_io_nasti_w_valid; // @[Tile.scala 128:19]
  wire [31:0] arb_io_nasti_w_bits_data; // @[Tile.scala 128:19]
  wire  arb_io_nasti_w_bits_last; // @[Tile.scala 128:19]
  wire  arb_io_nasti_b_ready; // @[Tile.scala 128:19]
  wire  arb_io_nasti_b_valid; // @[Tile.scala 128:19]
  wire  arb_io_nasti_ar_ready; // @[Tile.scala 128:19]
  wire  arb_io_nasti_ar_valid; // @[Tile.scala 128:19]
  wire [31:0] arb_io_nasti_ar_bits_addr; // @[Tile.scala 128:19]
  wire  arb_io_nasti_r_ready; // @[Tile.scala 128:19]
  wire  arb_io_nasti_r_valid; // @[Tile.scala 128:19]
  wire [31:0] arb_io_nasti_r_bits_data; // @[Tile.scala 128:19]
  wire  arb_io_nasti_r_bits_last; // @[Tile.scala 128:19]
  wire  selector_clock; // @[Tile.scala 129:24]
  wire  selector_reset; // @[Tile.scala 129:24]
  wire  selector_io_cpu_abort; // @[Tile.scala 129:24]
  wire  selector_io_cpu_req_valid; // @[Tile.scala 129:24]
  wire [31:0] selector_io_cpu_req_bits_addr; // @[Tile.scala 129:24]
  wire [31:0] selector_io_cpu_req_bits_data; // @[Tile.scala 129:24]
  wire [3:0] selector_io_cpu_req_bits_mask; // @[Tile.scala 129:24]
  wire  selector_io_cpu_resp_valid; // @[Tile.scala 129:24]
  wire [31:0] selector_io_cpu_resp_bits_data; // @[Tile.scala 129:24]
  wire  selector_io_dcache_abort; // @[Tile.scala 129:24]
  wire  selector_io_dcache_req_valid; // @[Tile.scala 129:24]
  wire [31:0] selector_io_dcache_req_bits_addr; // @[Tile.scala 129:24]
  wire [31:0] selector_io_dcache_req_bits_data; // @[Tile.scala 129:24]
  wire [3:0] selector_io_dcache_req_bits_mask; // @[Tile.scala 129:24]
  wire  selector_io_dcache_resp_valid; // @[Tile.scala 129:24]
  wire [31:0] selector_io_dcache_resp_bits_data; // @[Tile.scala 129:24]
  wire  selector_io_devices_req_valid; // @[Tile.scala 129:24]
  wire [31:0] selector_io_devices_req_bits_addr; // @[Tile.scala 129:24]
  wire [31:0] selector_io_devices_req_bits_data; // @[Tile.scala 129:24]
  wire [3:0] selector_io_devices_req_bits_mask; // @[Tile.scala 129:24]
  wire  selector_io_devices_resp_valid; // @[Tile.scala 129:24]
  wire [31:0] selector_io_devices_resp_bits_data; // @[Tile.scala 129:24]
  wire  immu_clock; // @[Tile.scala 130:20]
  wire  immu_reset; // @[Tile.scala 130:20]
  wire  immu_io_cpu_req_valid; // @[Tile.scala 130:20]
  wire [31:0] immu_io_cpu_req_bits_addr; // @[Tile.scala 130:20]
  wire  immu_io_cpu_resp_valid; // @[Tile.scala 130:20]
  wire [31:0] immu_io_cpu_resp_bits_data; // @[Tile.scala 130:20]
  wire  immu_io_cache_req_valid; // @[Tile.scala 130:20]
  wire [31:0] immu_io_cache_req_bits_addr; // @[Tile.scala 130:20]
  wire  immu_io_cache_resp_valid; // @[Tile.scala 130:20]
  wire [31:0] immu_io_cache_resp_bits_data; // @[Tile.scala 130:20]
  wire  immu_vmSwitch_0; // @[Tile.scala 130:20]
  wire [31:0] immu_csrWdata_0; // @[Tile.scala 130:20]
  wire  immu_clearPageFault_0; // @[Tile.scala 130:20]
  wire [1:0] immu_pageFault_1; // @[Tile.scala 130:20]
  wire [31:0] immu_satp_0; // @[Tile.scala 130:20]
  wire  dmmu_clock; // @[Tile.scala 131:20]
  wire  dmmu_reset; // @[Tile.scala 131:20]
  wire  dmmu_io_cpu_abort; // @[Tile.scala 131:20]
  wire  dmmu_io_cpu_req_valid; // @[Tile.scala 131:20]
  wire [31:0] dmmu_io_cpu_req_bits_addr; // @[Tile.scala 131:20]
  wire [31:0] dmmu_io_cpu_req_bits_data; // @[Tile.scala 131:20]
  wire [3:0] dmmu_io_cpu_req_bits_mask; // @[Tile.scala 131:20]
  wire  dmmu_io_cpu_resp_valid; // @[Tile.scala 131:20]
  wire [31:0] dmmu_io_cpu_resp_bits_data; // @[Tile.scala 131:20]
  wire  dmmu_io_cache_abort; // @[Tile.scala 131:20]
  wire  dmmu_io_cache_req_valid; // @[Tile.scala 131:20]
  wire [31:0] dmmu_io_cache_req_bits_addr; // @[Tile.scala 131:20]
  wire [31:0] dmmu_io_cache_req_bits_data; // @[Tile.scala 131:20]
  wire [3:0] dmmu_io_cache_req_bits_mask; // @[Tile.scala 131:20]
  wire  dmmu_io_cache_resp_valid; // @[Tile.scala 131:20]
  wire [31:0] dmmu_io_cache_resp_bits_data; // @[Tile.scala 131:20]
  wire [1:0] dmmu_pageFault_0; // @[Tile.scala 131:20]
  wire  dmmu_vmSwitch_0; // @[Tile.scala 131:20]
  wire [31:0] dmmu_csrWdata_0; // @[Tile.scala 131:20]
  wire  dmmu_clearPageFault_0; // @[Tile.scala 131:20]
  wire [31:0] dmmu_satp_0; // @[Tile.scala 131:20]
  wire  regmapper_clock; // @[Tile.scala 136:25]
  wire  regmapper_io_selector_req_valid; // @[Tile.scala 136:25]
  wire [31:0] regmapper_io_selector_req_bits_addr; // @[Tile.scala 136:25]
  wire [31:0] regmapper_io_selector_req_bits_data; // @[Tile.scala 136:25]
  wire [3:0] regmapper_io_selector_req_bits_mask; // @[Tile.scala 136:25]
  wire  regmapper_io_selector_resp_valid; // @[Tile.scala 136:25]
  wire [31:0] regmapper_io_selector_resp_bits_data; // @[Tile.scala 136:25]
  wire  regmapper_io_uart_req_valid; // @[Tile.scala 136:25]
  wire [31:0] regmapper_io_uart_req_bits_addr; // @[Tile.scala 136:25]
  wire [31:0] regmapper_io_uart_req_bits_data; // @[Tile.scala 136:25]
  wire  regmapper_io_uart_resp_valid; // @[Tile.scala 136:25]
  wire [31:0] regmapper_io_uart_resp_bits_data; // @[Tile.scala 136:25]
  wire  regmapper_io_rtc_req_valid; // @[Tile.scala 136:25]
  wire [31:0] regmapper_io_rtc_req_bits_addr; // @[Tile.scala 136:25]
  wire [31:0] regmapper_io_rtc_req_bits_data; // @[Tile.scala 136:25]
  wire [3:0] regmapper_io_rtc_req_bits_mask; // @[Tile.scala 136:25]
  wire  regmapper_io_rtc_resp_valid; // @[Tile.scala 136:25]
  wire [31:0] regmapper_io_rtc_resp_bits_data; // @[Tile.scala 136:25]
  wire  dram_io_nasti_aw_ready; // @[Tile.scala 139:20]
  wire  dram_io_nasti_aw_valid; // @[Tile.scala 139:20]
  wire [31:0] dram_io_nasti_aw_bits_addr; // @[Tile.scala 139:20]
  wire  dram_io_nasti_w_ready; // @[Tile.scala 139:20]
  wire  dram_io_nasti_w_valid; // @[Tile.scala 139:20]
  wire [31:0] dram_io_nasti_w_bits_data; // @[Tile.scala 139:20]
  wire  dram_io_nasti_w_bits_last; // @[Tile.scala 139:20]
  wire  dram_io_nasti_b_ready; // @[Tile.scala 139:20]
  wire  dram_io_nasti_b_valid; // @[Tile.scala 139:20]
  wire  dram_io_nasti_ar_ready; // @[Tile.scala 139:20]
  wire  dram_io_nasti_ar_valid; // @[Tile.scala 139:20]
  wire [31:0] dram_io_nasti_ar_bits_addr; // @[Tile.scala 139:20]
  wire  dram_io_nasti_r_ready; // @[Tile.scala 139:20]
  wire  dram_io_nasti_r_valid; // @[Tile.scala 139:20]
  wire [31:0] dram_io_nasti_r_bits_data; // @[Tile.scala 139:20]
  wire  dram_io_nasti_r_bits_last; // @[Tile.scala 139:20]
  wire [31:0] dram_io_AXI_s_axi_awaddr; // @[Tile.scala 139:20]
  wire  dram_io_AXI_s_axi_awvalid; // @[Tile.scala 139:20]
  wire  dram_io_AXI_s_axi_awready; // @[Tile.scala 139:20]
  wire [31:0] dram_io_AXI_s_axi_wdata; // @[Tile.scala 139:20]
  wire  dram_io_AXI_s_axi_wlast; // @[Tile.scala 139:20]
  wire  dram_io_AXI_s_axi_wvalid; // @[Tile.scala 139:20]
  wire  dram_io_AXI_s_axi_wready; // @[Tile.scala 139:20]
  wire  dram_io_AXI_s_axi_bvalid; // @[Tile.scala 139:20]
  wire  dram_io_AXI_s_axi_bready; // @[Tile.scala 139:20]
  wire [31:0] dram_io_AXI_s_axi_araddr; // @[Tile.scala 139:20]
  wire  dram_io_AXI_s_axi_arvalid; // @[Tile.scala 139:20]
  wire  dram_io_AXI_s_axi_arready; // @[Tile.scala 139:20]
  wire [31:0] dram_io_AXI_s_axi_rdata; // @[Tile.scala 139:20]
  wire  dram_io_AXI_s_axi_rlast; // @[Tile.scala 139:20]
  wire  dram_io_AXI_s_axi_rvalid; // @[Tile.scala 139:20]
  wire  dram_io_AXI_s_axi_rready; // @[Tile.scala 139:20]
  wire  uartController_clock; // @[Tile.scala 142:30]
  wire  uartController_reset; // @[Tile.scala 142:30]
  wire  uartController_io__cpu_req_valid; // @[Tile.scala 142:30]
  wire [31:0] uartController_io__cpu_req_bits_addr; // @[Tile.scala 142:30]
  wire [31:0] uartController_io__cpu_req_bits_data; // @[Tile.scala 142:30]
  wire  uartController_io__cpu_resp_valid; // @[Tile.scala 142:30]
  wire [31:0] uartController_io__cpu_resp_bits_data; // @[Tile.scala 142:30]
  wire  uartController_io__rxChannel_ready; // @[Tile.scala 142:30]
  wire  uartController_io__rxChannel_valid; // @[Tile.scala 142:30]
  wire [7:0] uartController_io__rxChannel_bits; // @[Tile.scala 142:30]
  wire  uartController_io__txChannel_ready; // @[Tile.scala 142:30]
  wire  uartController_io__txChannel_valid; // @[Tile.scala 142:30]
  wire [7:0] uartController_io__txChannel_bits; // @[Tile.scala 142:30]
  wire  uartController_io_rxChannel_valid; // @[Tile.scala 142:30]
  wire  uart_clock; // @[Tile.scala 143:20]
  wire  uart_reset; // @[Tile.scala 143:20]
  wire  uart_io_rxd; // @[Tile.scala 143:20]
  wire  uart_io_txd; // @[Tile.scala 143:20]
  wire  uart_io_rxChannel_ready; // @[Tile.scala 143:20]
  wire  uart_io_rxChannel_valid; // @[Tile.scala 143:20]
  wire [7:0] uart_io_rxChannel_bits; // @[Tile.scala 143:20]
  wire  uart_io_txChannel_ready; // @[Tile.scala 143:20]
  wire  uart_io_txChannel_valid; // @[Tile.scala 143:20]
  wire [7:0] uart_io_txChannel_bits; // @[Tile.scala 143:20]
  wire  rtc_clock; // @[Tile.scala 145:19]
  wire  rtc_reset; // @[Tile.scala 145:19]
  wire  rtc_io_req_valid; // @[Tile.scala 145:19]
  wire [31:0] rtc_io_req_bits_addr; // @[Tile.scala 145:19]
  wire [31:0] rtc_io_req_bits_data; // @[Tile.scala 145:19]
  wire [3:0] rtc_io_req_bits_mask; // @[Tile.scala 145:19]
  wire  rtc_io_resp_valid; // @[Tile.scala 145:19]
  wire [31:0] rtc_io_resp_bits_data; // @[Tile.scala 145:19]
  DFC_Table dfc_table ( // @[Tile.scala 120:25]
    .clock(dfc_table_clock),
    .reset(dfc_table_reset),
    .io_cpu1_w_data_valid(dfc_table_io_cpu1_w_data_valid),
    .io_cpu1_w_data_bits_listenAddr(dfc_table_io_cpu1_w_data_bits_listenAddr),
    .io_cpu1_w_data_bits_wPid(dfc_table_io_cpu1_w_data_bits_wPid),
    .io_cpu1_l_data_valid(dfc_table_io_cpu1_l_data_valid),
    .io_cpu1_l_data_bits_listenAddr(dfc_table_io_cpu1_l_data_bits_listenAddr),
    .io_cpu1_e_data_ready(dfc_table_io_cpu1_e_data_ready),
    .io_cpu1_e_data_valid(dfc_table_io_cpu1_e_data_valid),
    .io_cpu1_e_data_bits_pid(dfc_table_io_cpu1_e_data_bits_pid),
    .io_cpu_f_data_valid(dfc_table_io_cpu_f_data_valid),
    .io_cpu_f_data_bits_full_sig(dfc_table_io_cpu_f_data_bits_full_sig)
  );
  Core core ( // @[Tile.scala 125:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_icache_req_valid(core_io_icache_req_valid),
    .io_icache_req_bits_addr(core_io_icache_req_bits_addr),
    .io_icache_resp_valid(core_io_icache_resp_valid),
    .io_icache_resp_bits_data(core_io_icache_resp_bits_data),
    .io_dcache_abort(core_io_dcache_abort),
    .io_dcache_req_valid(core_io_dcache_req_valid),
    .io_dcache_req_bits_addr(core_io_dcache_req_bits_addr),
    .io_dcache_req_bits_data(core_io_dcache_req_bits_data),
    .io_dcache_req_bits_mask(core_io_dcache_req_bits_mask),
    .io_dcache_resp_valid(core_io_dcache_resp_valid),
    .io_dcache_resp_bits_data(core_io_dcache_resp_bits_data),
    .io_table_w_data_valid(core_io_table_w_data_valid),
    .io_table_w_data_bits_listenAddr(core_io_table_w_data_bits_listenAddr),
    .io_table_w_data_bits_wPid(core_io_table_w_data_bits_wPid),
    .io_table_l_data_valid(core_io_table_l_data_valid),
    .io_table_l_data_bits_listenAddr(core_io_table_l_data_bits_listenAddr),
    .io_table_e_data_ready(core_io_table_e_data_ready),
    .io_table_e_data_valid(core_io_table_e_data_valid),
    .io_table_e_data_bits_pid(core_io_table_e_data_bits_pid),
    .io_table_f_data_valid(core_io_table_f_data_valid),
    .io_table_f_data_bits_full_sig(core_io_table_f_data_bits_full_sig),
    .io_rxChannel_valid(core_io_rxChannel_valid),
    .pageFault(core_pageFault),
    .io_vmSwitch(core_io_vmSwitch),
    .io_in(core_io_in),
    .clearPageFault(core_clearPageFault),
    .pageFault_0(core_pageFault_0),
    .satp(core_satp)
  );
  Cache icache ( // @[Tile.scala 126:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_cpu_abort(icache_io_cpu_abort),
    .io_cpu_req_valid(icache_io_cpu_req_valid),
    .io_cpu_req_bits_addr(icache_io_cpu_req_bits_addr),
    .io_cpu_req_bits_data(icache_io_cpu_req_bits_data),
    .io_cpu_req_bits_mask(icache_io_cpu_req_bits_mask),
    .io_cpu_resp_valid(icache_io_cpu_resp_valid),
    .io_cpu_resp_bits_data(icache_io_cpu_resp_bits_data),
    .io_nasti_aw_ready(icache_io_nasti_aw_ready),
    .io_nasti_aw_valid(icache_io_nasti_aw_valid),
    .io_nasti_aw_bits_addr(icache_io_nasti_aw_bits_addr),
    .io_nasti_w_ready(icache_io_nasti_w_ready),
    .io_nasti_w_valid(icache_io_nasti_w_valid),
    .io_nasti_w_bits_data(icache_io_nasti_w_bits_data),
    .io_nasti_w_bits_last(icache_io_nasti_w_bits_last),
    .io_nasti_b_ready(icache_io_nasti_b_ready),
    .io_nasti_b_valid(icache_io_nasti_b_valid),
    .io_nasti_ar_ready(icache_io_nasti_ar_ready),
    .io_nasti_ar_valid(icache_io_nasti_ar_valid),
    .io_nasti_ar_bits_addr(icache_io_nasti_ar_bits_addr),
    .io_nasti_r_ready(icache_io_nasti_r_ready),
    .io_nasti_r_valid(icache_io_nasti_r_valid),
    .io_nasti_r_bits_data(icache_io_nasti_r_bits_data)
  );
  Cache dcache ( // @[Tile.scala 127:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_cpu_abort(dcache_io_cpu_abort),
    .io_cpu_req_valid(dcache_io_cpu_req_valid),
    .io_cpu_req_bits_addr(dcache_io_cpu_req_bits_addr),
    .io_cpu_req_bits_data(dcache_io_cpu_req_bits_data),
    .io_cpu_req_bits_mask(dcache_io_cpu_req_bits_mask),
    .io_cpu_resp_valid(dcache_io_cpu_resp_valid),
    .io_cpu_resp_bits_data(dcache_io_cpu_resp_bits_data),
    .io_nasti_aw_ready(dcache_io_nasti_aw_ready),
    .io_nasti_aw_valid(dcache_io_nasti_aw_valid),
    .io_nasti_aw_bits_addr(dcache_io_nasti_aw_bits_addr),
    .io_nasti_w_ready(dcache_io_nasti_w_ready),
    .io_nasti_w_valid(dcache_io_nasti_w_valid),
    .io_nasti_w_bits_data(dcache_io_nasti_w_bits_data),
    .io_nasti_w_bits_last(dcache_io_nasti_w_bits_last),
    .io_nasti_b_ready(dcache_io_nasti_b_ready),
    .io_nasti_b_valid(dcache_io_nasti_b_valid),
    .io_nasti_ar_ready(dcache_io_nasti_ar_ready),
    .io_nasti_ar_valid(dcache_io_nasti_ar_valid),
    .io_nasti_ar_bits_addr(dcache_io_nasti_ar_bits_addr),
    .io_nasti_r_ready(dcache_io_nasti_r_ready),
    .io_nasti_r_valid(dcache_io_nasti_r_valid),
    .io_nasti_r_bits_data(dcache_io_nasti_r_bits_data)
  );
  MemArbiter arb ( // @[Tile.scala 128:19]
    .clock(arb_clock),
    .reset(arb_reset),
    .io_icache_ar_ready(arb_io_icache_ar_ready),
    .io_icache_ar_valid(arb_io_icache_ar_valid),
    .io_icache_ar_bits_addr(arb_io_icache_ar_bits_addr),
    .io_icache_r_ready(arb_io_icache_r_ready),
    .io_icache_r_valid(arb_io_icache_r_valid),
    .io_icache_r_bits_data(arb_io_icache_r_bits_data),
    .io_dcache_aw_ready(arb_io_dcache_aw_ready),
    .io_dcache_aw_valid(arb_io_dcache_aw_valid),
    .io_dcache_aw_bits_addr(arb_io_dcache_aw_bits_addr),
    .io_dcache_w_ready(arb_io_dcache_w_ready),
    .io_dcache_w_valid(arb_io_dcache_w_valid),
    .io_dcache_w_bits_data(arb_io_dcache_w_bits_data),
    .io_dcache_w_bits_last(arb_io_dcache_w_bits_last),
    .io_dcache_b_ready(arb_io_dcache_b_ready),
    .io_dcache_b_valid(arb_io_dcache_b_valid),
    .io_dcache_ar_ready(arb_io_dcache_ar_ready),
    .io_dcache_ar_valid(arb_io_dcache_ar_valid),
    .io_dcache_ar_bits_addr(arb_io_dcache_ar_bits_addr),
    .io_dcache_r_ready(arb_io_dcache_r_ready),
    .io_dcache_r_valid(arb_io_dcache_r_valid),
    .io_dcache_r_bits_data(arb_io_dcache_r_bits_data),
    .io_nasti_aw_ready(arb_io_nasti_aw_ready),
    .io_nasti_aw_valid(arb_io_nasti_aw_valid),
    .io_nasti_aw_bits_addr(arb_io_nasti_aw_bits_addr),
    .io_nasti_w_ready(arb_io_nasti_w_ready),
    .io_nasti_w_valid(arb_io_nasti_w_valid),
    .io_nasti_w_bits_data(arb_io_nasti_w_bits_data),
    .io_nasti_w_bits_last(arb_io_nasti_w_bits_last),
    .io_nasti_b_ready(arb_io_nasti_b_ready),
    .io_nasti_b_valid(arb_io_nasti_b_valid),
    .io_nasti_ar_ready(arb_io_nasti_ar_ready),
    .io_nasti_ar_valid(arb_io_nasti_ar_valid),
    .io_nasti_ar_bits_addr(arb_io_nasti_ar_bits_addr),
    .io_nasti_r_ready(arb_io_nasti_r_ready),
    .io_nasti_r_valid(arb_io_nasti_r_valid),
    .io_nasti_r_bits_data(arb_io_nasti_r_bits_data),
    .io_nasti_r_bits_last(arb_io_nasti_r_bits_last)
  );
  Selector selector ( // @[Tile.scala 129:24]
    .clock(selector_clock),
    .reset(selector_reset),
    .io_cpu_abort(selector_io_cpu_abort),
    .io_cpu_req_valid(selector_io_cpu_req_valid),
    .io_cpu_req_bits_addr(selector_io_cpu_req_bits_addr),
    .io_cpu_req_bits_data(selector_io_cpu_req_bits_data),
    .io_cpu_req_bits_mask(selector_io_cpu_req_bits_mask),
    .io_cpu_resp_valid(selector_io_cpu_resp_valid),
    .io_cpu_resp_bits_data(selector_io_cpu_resp_bits_data),
    .io_dcache_abort(selector_io_dcache_abort),
    .io_dcache_req_valid(selector_io_dcache_req_valid),
    .io_dcache_req_bits_addr(selector_io_dcache_req_bits_addr),
    .io_dcache_req_bits_data(selector_io_dcache_req_bits_data),
    .io_dcache_req_bits_mask(selector_io_dcache_req_bits_mask),
    .io_dcache_resp_valid(selector_io_dcache_resp_valid),
    .io_dcache_resp_bits_data(selector_io_dcache_resp_bits_data),
    .io_devices_req_valid(selector_io_devices_req_valid),
    .io_devices_req_bits_addr(selector_io_devices_req_bits_addr),
    .io_devices_req_bits_data(selector_io_devices_req_bits_data),
    .io_devices_req_bits_mask(selector_io_devices_req_bits_mask),
    .io_devices_resp_valid(selector_io_devices_resp_valid),
    .io_devices_resp_bits_data(selector_io_devices_resp_bits_data)
  );
  MMU immu ( // @[Tile.scala 130:20]
    .clock(immu_clock),
    .reset(immu_reset),
    .io_cpu_req_valid(immu_io_cpu_req_valid),
    .io_cpu_req_bits_addr(immu_io_cpu_req_bits_addr),
    .io_cpu_resp_valid(immu_io_cpu_resp_valid),
    .io_cpu_resp_bits_data(immu_io_cpu_resp_bits_data),
    .io_cache_req_valid(immu_io_cache_req_valid),
    .io_cache_req_bits_addr(immu_io_cache_req_bits_addr),
    .io_cache_resp_valid(immu_io_cache_resp_valid),
    .io_cache_resp_bits_data(immu_io_cache_resp_bits_data),
    .vmSwitch_0(immu_vmSwitch_0),
    .csrWdata_0(immu_csrWdata_0),
    .clearPageFault_0(immu_clearPageFault_0),
    .pageFault_1(immu_pageFault_1),
    .satp_0(immu_satp_0)
  );
  MMU_1 dmmu ( // @[Tile.scala 131:20]
    .clock(dmmu_clock),
    .reset(dmmu_reset),
    .io_cpu_abort(dmmu_io_cpu_abort),
    .io_cpu_req_valid(dmmu_io_cpu_req_valid),
    .io_cpu_req_bits_addr(dmmu_io_cpu_req_bits_addr),
    .io_cpu_req_bits_data(dmmu_io_cpu_req_bits_data),
    .io_cpu_req_bits_mask(dmmu_io_cpu_req_bits_mask),
    .io_cpu_resp_valid(dmmu_io_cpu_resp_valid),
    .io_cpu_resp_bits_data(dmmu_io_cpu_resp_bits_data),
    .io_cache_abort(dmmu_io_cache_abort),
    .io_cache_req_valid(dmmu_io_cache_req_valid),
    .io_cache_req_bits_addr(dmmu_io_cache_req_bits_addr),
    .io_cache_req_bits_data(dmmu_io_cache_req_bits_data),
    .io_cache_req_bits_mask(dmmu_io_cache_req_bits_mask),
    .io_cache_resp_valid(dmmu_io_cache_resp_valid),
    .io_cache_resp_bits_data(dmmu_io_cache_resp_bits_data),
    .pageFault_0(dmmu_pageFault_0),
    .vmSwitch_0(dmmu_vmSwitch_0),
    .csrWdata_0(dmmu_csrWdata_0),
    .clearPageFault_0(dmmu_clearPageFault_0),
    .satp_0(dmmu_satp_0)
  );
  RegMapper regmapper ( // @[Tile.scala 136:25]
    .clock(regmapper_clock),
    .io_selector_req_valid(regmapper_io_selector_req_valid),
    .io_selector_req_bits_addr(regmapper_io_selector_req_bits_addr),
    .io_selector_req_bits_data(regmapper_io_selector_req_bits_data),
    .io_selector_req_bits_mask(regmapper_io_selector_req_bits_mask),
    .io_selector_resp_valid(regmapper_io_selector_resp_valid),
    .io_selector_resp_bits_data(regmapper_io_selector_resp_bits_data),
    .io_uart_req_valid(regmapper_io_uart_req_valid),
    .io_uart_req_bits_addr(regmapper_io_uart_req_bits_addr),
    .io_uart_req_bits_data(regmapper_io_uart_req_bits_data),
    .io_uart_resp_valid(regmapper_io_uart_resp_valid),
    .io_uart_resp_bits_data(regmapper_io_uart_resp_bits_data),
    .io_rtc_req_valid(regmapper_io_rtc_req_valid),
    .io_rtc_req_bits_addr(regmapper_io_rtc_req_bits_addr),
    .io_rtc_req_bits_data(regmapper_io_rtc_req_bits_data),
    .io_rtc_req_bits_mask(regmapper_io_rtc_req_bits_mask),
    .io_rtc_resp_valid(regmapper_io_rtc_resp_valid),
    .io_rtc_resp_bits_data(regmapper_io_rtc_resp_bits_data)
  );
  DRAM dram ( // @[Tile.scala 139:20]
    .io_nasti_aw_ready(dram_io_nasti_aw_ready),
    .io_nasti_aw_valid(dram_io_nasti_aw_valid),
    .io_nasti_aw_bits_addr(dram_io_nasti_aw_bits_addr),
    .io_nasti_w_ready(dram_io_nasti_w_ready),
    .io_nasti_w_valid(dram_io_nasti_w_valid),
    .io_nasti_w_bits_data(dram_io_nasti_w_bits_data),
    .io_nasti_w_bits_last(dram_io_nasti_w_bits_last),
    .io_nasti_b_ready(dram_io_nasti_b_ready),
    .io_nasti_b_valid(dram_io_nasti_b_valid),
    .io_nasti_ar_ready(dram_io_nasti_ar_ready),
    .io_nasti_ar_valid(dram_io_nasti_ar_valid),
    .io_nasti_ar_bits_addr(dram_io_nasti_ar_bits_addr),
    .io_nasti_r_ready(dram_io_nasti_r_ready),
    .io_nasti_r_valid(dram_io_nasti_r_valid),
    .io_nasti_r_bits_data(dram_io_nasti_r_bits_data),
    .io_nasti_r_bits_last(dram_io_nasti_r_bits_last),
    .io_AXI_s_axi_awaddr(dram_io_AXI_s_axi_awaddr),
    .io_AXI_s_axi_awvalid(dram_io_AXI_s_axi_awvalid),
    .io_AXI_s_axi_awready(dram_io_AXI_s_axi_awready),
    .io_AXI_s_axi_wdata(dram_io_AXI_s_axi_wdata),
    .io_AXI_s_axi_wlast(dram_io_AXI_s_axi_wlast),
    .io_AXI_s_axi_wvalid(dram_io_AXI_s_axi_wvalid),
    .io_AXI_s_axi_wready(dram_io_AXI_s_axi_wready),
    .io_AXI_s_axi_bvalid(dram_io_AXI_s_axi_bvalid),
    .io_AXI_s_axi_bready(dram_io_AXI_s_axi_bready),
    .io_AXI_s_axi_araddr(dram_io_AXI_s_axi_araddr),
    .io_AXI_s_axi_arvalid(dram_io_AXI_s_axi_arvalid),
    .io_AXI_s_axi_arready(dram_io_AXI_s_axi_arready),
    .io_AXI_s_axi_rdata(dram_io_AXI_s_axi_rdata),
    .io_AXI_s_axi_rlast(dram_io_AXI_s_axi_rlast),
    .io_AXI_s_axi_rvalid(dram_io_AXI_s_axi_rvalid),
    .io_AXI_s_axi_rready(dram_io_AXI_s_axi_rready)
  );
  UartController uartController ( // @[Tile.scala 142:30]
    .clock(uartController_clock),
    .reset(uartController_reset),
    .io__cpu_req_valid(uartController_io__cpu_req_valid),
    .io__cpu_req_bits_addr(uartController_io__cpu_req_bits_addr),
    .io__cpu_req_bits_data(uartController_io__cpu_req_bits_data),
    .io__cpu_resp_valid(uartController_io__cpu_resp_valid),
    .io__cpu_resp_bits_data(uartController_io__cpu_resp_bits_data),
    .io__rxChannel_ready(uartController_io__rxChannel_ready),
    .io__rxChannel_valid(uartController_io__rxChannel_valid),
    .io__rxChannel_bits(uartController_io__rxChannel_bits),
    .io__txChannel_ready(uartController_io__txChannel_ready),
    .io__txChannel_valid(uartController_io__txChannel_valid),
    .io__txChannel_bits(uartController_io__txChannel_bits),
    .io_rxChannel_valid(uartController_io_rxChannel_valid)
  );
  Uart uart ( // @[Tile.scala 143:20]
    .clock(uart_clock),
    .reset(uart_reset),
    .io_rxd(uart_io_rxd),
    .io_txd(uart_io_txd),
    .io_rxChannel_ready(uart_io_rxChannel_ready),
    .io_rxChannel_valid(uart_io_rxChannel_valid),
    .io_rxChannel_bits(uart_io_rxChannel_bits),
    .io_txChannel_ready(uart_io_txChannel_ready),
    .io_txChannel_valid(uart_io_txChannel_valid),
    .io_txChannel_bits(uart_io_txChannel_bits)
  );
  RTC rtc ( // @[Tile.scala 145:19]
    .clock(rtc_clock),
    .reset(rtc_reset),
    .io_req_valid(rtc_io_req_valid),
    .io_req_bits_addr(rtc_io_req_bits_addr),
    .io_req_bits_data(rtc_io_req_bits_data),
    .io_req_bits_mask(rtc_io_req_bits_mask),
    .io_resp_valid(rtc_io_resp_valid),
    .io_resp_bits_data(rtc_io_resp_bits_data)
  );
  assign io_AXI_s_axi_awid = 4'h0; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_awaddr = dram_io_AXI_s_axi_awaddr; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_awlen = 8'h0; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_awsize = 3'h2; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_awburst = 2'h1; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_awvalid = dram_io_AXI_s_axi_awvalid; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_wdata = dram_io_AXI_s_axi_wdata; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_wstrb = 8'hf; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_wlast = dram_io_AXI_s_axi_wlast; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_wvalid = dram_io_AXI_s_axi_wvalid; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_bready = dram_io_AXI_s_axi_bready; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_arid = 4'h0; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_araddr = dram_io_AXI_s_axi_araddr; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_arlen = 8'h0; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_arsize = 3'h2; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_arburst = 2'h1; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_arvalid = dram_io_AXI_s_axi_arvalid; // @[Tile.scala 187:10]
  assign io_AXI_s_axi_rready = dram_io_AXI_s_axi_rready; // @[Tile.scala 187:10]
  assign io_txd = uart_io_txd; // @[Tile.scala 173:15]
  assign dfc_table_clock = clock;
  assign dfc_table_reset = reset;
  assign dfc_table_io_cpu1_w_data_valid = core_io_table_w_data_valid; // @[Tile.scala 190:23]
  assign dfc_table_io_cpu1_w_data_bits_listenAddr = core_io_table_w_data_bits_listenAddr; // @[Tile.scala 190:23]
  assign dfc_table_io_cpu1_w_data_bits_wPid = core_io_table_w_data_bits_wPid; // @[Tile.scala 190:23]
  assign dfc_table_io_cpu1_l_data_valid = core_io_table_l_data_valid; // @[Tile.scala 191:23]
  assign dfc_table_io_cpu1_l_data_bits_listenAddr = core_io_table_l_data_bits_listenAddr; // @[Tile.scala 191:23]
  assign dfc_table_io_cpu1_e_data_ready = core_io_table_e_data_ready; // @[Tile.scala 201:19]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_icache_resp_valid = immu_io_cpu_resp_valid; // @[Tile.scala 158:18]
  assign core_io_icache_resp_bits_data = immu_io_cpu_resp_bits_data; // @[Tile.scala 158:18]
  assign core_io_dcache_resp_valid = selector_io_cpu_resp_valid; // @[Tile.scala 160:18]
  assign core_io_dcache_resp_bits_data = selector_io_cpu_resp_bits_data; // @[Tile.scala 160:18]
  assign core_io_table_e_data_valid = dfc_table_io_cpu1_e_data_valid; // @[Tile.scala 201:19]
  assign core_io_table_e_data_bits_pid = dfc_table_io_cpu1_e_data_bits_pid; // @[Tile.scala 201:19]
  assign core_io_table_f_data_valid = dfc_table_io_cpu_f_data_valid; // @[Tile.scala 202:19]
  assign core_io_table_f_data_bits_full_sig = dfc_table_io_cpu_f_data_bits_full_sig; // @[Tile.scala 202:19]
  assign core_io_rxChannel_valid = uartController_io_rxChannel_valid;
  assign core_pageFault = dmmu_pageFault_0;
  assign core_pageFault_0 = immu_pageFault_1;
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_cpu_abort = 1'h0; // @[Tile.scala 159:17]
  assign icache_io_cpu_req_valid = immu_io_cache_req_valid; // @[Tile.scala 159:17]
  assign icache_io_cpu_req_bits_addr = immu_io_cache_req_bits_addr; // @[Tile.scala 159:17]
  assign icache_io_cpu_req_bits_data = 32'h0; // @[Tile.scala 159:17]
  assign icache_io_cpu_req_bits_mask = 4'h0; // @[Tile.scala 159:17]
  assign icache_io_nasti_aw_ready = 1'h0; // @[Tile.scala 180:17]
  assign icache_io_nasti_w_ready = 1'h0; // @[Tile.scala 180:17]
  assign icache_io_nasti_b_valid = 1'h0; // @[Tile.scala 180:17]
  assign icache_io_nasti_ar_ready = arb_io_icache_ar_ready; // @[Tile.scala 180:17]
  assign icache_io_nasti_r_valid = arb_io_icache_r_valid; // @[Tile.scala 180:17]
  assign icache_io_nasti_r_bits_data = arb_io_icache_r_bits_data; // @[Tile.scala 180:17]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_cpu_abort = dmmu_io_cache_abort; // @[Tile.scala 165:17]
  assign dcache_io_cpu_req_valid = dmmu_io_cache_req_valid; // @[Tile.scala 165:17]
  assign dcache_io_cpu_req_bits_addr = dmmu_io_cache_req_bits_addr; // @[Tile.scala 165:17]
  assign dcache_io_cpu_req_bits_data = dmmu_io_cache_req_bits_data; // @[Tile.scala 165:17]
  assign dcache_io_cpu_req_bits_mask = dmmu_io_cache_req_bits_mask; // @[Tile.scala 165:17]
  assign dcache_io_nasti_aw_ready = arb_io_dcache_aw_ready; // @[Tile.scala 181:17]
  assign dcache_io_nasti_w_ready = arb_io_dcache_w_ready; // @[Tile.scala 181:17]
  assign dcache_io_nasti_b_valid = arb_io_dcache_b_valid; // @[Tile.scala 181:17]
  assign dcache_io_nasti_ar_ready = arb_io_dcache_ar_ready; // @[Tile.scala 181:17]
  assign dcache_io_nasti_r_valid = arb_io_dcache_r_valid; // @[Tile.scala 181:17]
  assign dcache_io_nasti_r_bits_data = arb_io_dcache_r_bits_data; // @[Tile.scala 181:17]
  assign arb_clock = clock;
  assign arb_reset = reset;
  assign arb_io_icache_ar_valid = icache_io_nasti_ar_valid; // @[Tile.scala 180:17]
  assign arb_io_icache_ar_bits_addr = icache_io_nasti_ar_bits_addr; // @[Tile.scala 180:17]
  assign arb_io_icache_r_ready = icache_io_nasti_r_ready; // @[Tile.scala 180:17]
  assign arb_io_dcache_aw_valid = dcache_io_nasti_aw_valid; // @[Tile.scala 181:17]
  assign arb_io_dcache_aw_bits_addr = dcache_io_nasti_aw_bits_addr; // @[Tile.scala 181:17]
  assign arb_io_dcache_w_valid = dcache_io_nasti_w_valid; // @[Tile.scala 181:17]
  assign arb_io_dcache_w_bits_data = dcache_io_nasti_w_bits_data; // @[Tile.scala 181:17]
  assign arb_io_dcache_w_bits_last = dcache_io_nasti_w_bits_last; // @[Tile.scala 181:17]
  assign arb_io_dcache_b_ready = dcache_io_nasti_b_ready; // @[Tile.scala 181:17]
  assign arb_io_dcache_ar_valid = dcache_io_nasti_ar_valid; // @[Tile.scala 181:17]
  assign arb_io_dcache_ar_bits_addr = dcache_io_nasti_ar_bits_addr; // @[Tile.scala 181:17]
  assign arb_io_dcache_r_ready = dcache_io_nasti_r_ready; // @[Tile.scala 181:17]
  assign arb_io_nasti_aw_ready = dram_io_nasti_aw_ready; // @[Tile.scala 186:17]
  assign arb_io_nasti_w_ready = dram_io_nasti_w_ready; // @[Tile.scala 186:17]
  assign arb_io_nasti_b_valid = dram_io_nasti_b_valid; // @[Tile.scala 186:17]
  assign arb_io_nasti_ar_ready = dram_io_nasti_ar_ready; // @[Tile.scala 186:17]
  assign arb_io_nasti_r_valid = dram_io_nasti_r_valid; // @[Tile.scala 186:17]
  assign arb_io_nasti_r_bits_data = dram_io_nasti_r_bits_data; // @[Tile.scala 186:17]
  assign arb_io_nasti_r_bits_last = dram_io_nasti_r_bits_last; // @[Tile.scala 186:17]
  assign selector_clock = clock;
  assign selector_reset = reset;
  assign selector_io_cpu_abort = core_io_dcache_abort; // @[Tile.scala 160:18]
  assign selector_io_cpu_req_valid = core_io_dcache_req_valid; // @[Tile.scala 160:18]
  assign selector_io_cpu_req_bits_addr = core_io_dcache_req_bits_addr; // @[Tile.scala 160:18]
  assign selector_io_cpu_req_bits_data = core_io_dcache_req_bits_data; // @[Tile.scala 160:18]
  assign selector_io_cpu_req_bits_mask = core_io_dcache_req_bits_mask; // @[Tile.scala 160:18]
  assign selector_io_dcache_resp_valid = dmmu_io_cpu_resp_valid; // @[Tile.scala 164:22]
  assign selector_io_dcache_resp_bits_data = dmmu_io_cpu_resp_bits_data; // @[Tile.scala 164:22]
  assign selector_io_devices_resp_valid = regmapper_io_selector_resp_valid; // @[Tile.scala 166:23]
  assign selector_io_devices_resp_bits_data = regmapper_io_selector_resp_bits_data; // @[Tile.scala 166:23]
  assign immu_clock = clock;
  assign immu_reset = reset;
  assign immu_io_cpu_req_valid = core_io_icache_req_valid; // @[Tile.scala 158:18]
  assign immu_io_cpu_req_bits_addr = core_io_icache_req_bits_addr; // @[Tile.scala 158:18]
  assign immu_io_cache_resp_valid = icache_io_cpu_resp_valid; // @[Tile.scala 159:17]
  assign immu_io_cache_resp_bits_data = icache_io_cpu_resp_bits_data; // @[Tile.scala 159:17]
  assign immu_vmSwitch_0 = core_io_vmSwitch;
  assign immu_csrWdata_0 = core_io_in;
  assign immu_clearPageFault_0 = core_clearPageFault;
  assign immu_satp_0 = core_satp;
  assign dmmu_clock = clock;
  assign dmmu_reset = reset;
  assign dmmu_io_cpu_abort = selector_io_dcache_abort; // @[Tile.scala 164:22]
  assign dmmu_io_cpu_req_valid = selector_io_dcache_req_valid; // @[Tile.scala 164:22]
  assign dmmu_io_cpu_req_bits_addr = selector_io_dcache_req_bits_addr; // @[Tile.scala 164:22]
  assign dmmu_io_cpu_req_bits_data = selector_io_dcache_req_bits_data; // @[Tile.scala 164:22]
  assign dmmu_io_cpu_req_bits_mask = selector_io_dcache_req_bits_mask; // @[Tile.scala 164:22]
  assign dmmu_io_cache_resp_valid = dcache_io_cpu_resp_valid; // @[Tile.scala 165:17]
  assign dmmu_io_cache_resp_bits_data = dcache_io_cpu_resp_bits_data; // @[Tile.scala 165:17]
  assign dmmu_vmSwitch_0 = core_io_vmSwitch;
  assign dmmu_csrWdata_0 = core_io_in;
  assign dmmu_clearPageFault_0 = core_clearPageFault;
  assign dmmu_satp_0 = core_satp;
  assign regmapper_clock = clock;
  assign regmapper_io_selector_req_valid = selector_io_devices_req_valid; // @[Tile.scala 166:23]
  assign regmapper_io_selector_req_bits_addr = selector_io_devices_req_bits_addr; // @[Tile.scala 166:23]
  assign regmapper_io_selector_req_bits_data = selector_io_devices_req_bits_data; // @[Tile.scala 166:23]
  assign regmapper_io_selector_req_bits_mask = selector_io_devices_req_bits_mask; // @[Tile.scala 166:23]
  assign regmapper_io_uart_resp_valid = uartController_io__cpu_resp_valid; // @[Tile.scala 168:21]
  assign regmapper_io_uart_resp_bits_data = uartController_io__cpu_resp_bits_data; // @[Tile.scala 168:21]
  assign regmapper_io_rtc_resp_valid = rtc_io_resp_valid; // @[Tile.scala 177:20]
  assign regmapper_io_rtc_resp_bits_data = rtc_io_resp_bits_data; // @[Tile.scala 177:20]
  assign dram_io_nasti_aw_valid = arb_io_nasti_aw_valid; // @[Tile.scala 186:17]
  assign dram_io_nasti_aw_bits_addr = arb_io_nasti_aw_bits_addr; // @[Tile.scala 186:17]
  assign dram_io_nasti_w_valid = arb_io_nasti_w_valid; // @[Tile.scala 186:17]
  assign dram_io_nasti_w_bits_data = arb_io_nasti_w_bits_data; // @[Tile.scala 186:17]
  assign dram_io_nasti_w_bits_last = arb_io_nasti_w_bits_last; // @[Tile.scala 186:17]
  assign dram_io_nasti_b_ready = arb_io_nasti_b_ready; // @[Tile.scala 186:17]
  assign dram_io_nasti_ar_valid = arb_io_nasti_ar_valid; // @[Tile.scala 186:17]
  assign dram_io_nasti_ar_bits_addr = arb_io_nasti_ar_bits_addr; // @[Tile.scala 186:17]
  assign dram_io_nasti_r_ready = arb_io_nasti_r_ready; // @[Tile.scala 186:17]
  assign dram_io_AXI_s_axi_awready = io_AXI_s_axi_awready; // @[Tile.scala 187:10]
  assign dram_io_AXI_s_axi_wready = io_AXI_s_axi_wready; // @[Tile.scala 187:10]
  assign dram_io_AXI_s_axi_bvalid = io_AXI_s_axi_bvalid; // @[Tile.scala 187:10]
  assign dram_io_AXI_s_axi_arready = io_AXI_s_axi_arready; // @[Tile.scala 187:10]
  assign dram_io_AXI_s_axi_rdata = io_AXI_s_axi_rdata; // @[Tile.scala 187:10]
  assign dram_io_AXI_s_axi_rlast = io_AXI_s_axi_rlast; // @[Tile.scala 187:10]
  assign dram_io_AXI_s_axi_rvalid = io_AXI_s_axi_rvalid; // @[Tile.scala 187:10]
  assign uartController_clock = clock;
  assign uartController_reset = reset;
  assign uartController_io__cpu_req_valid = regmapper_io_uart_req_valid; // @[Tile.scala 168:21]
  assign uartController_io__cpu_req_bits_addr = regmapper_io_uart_req_bits_addr; // @[Tile.scala 168:21]
  assign uartController_io__cpu_req_bits_data = regmapper_io_uart_req_bits_data; // @[Tile.scala 168:21]
  assign uartController_io__rxChannel_valid = uart_io_rxChannel_valid; // @[Tile.scala 170:31]
  assign uartController_io__rxChannel_bits = uart_io_rxChannel_bits; // @[Tile.scala 170:31]
  assign uartController_io__txChannel_ready = uart_io_txChannel_ready; // @[Tile.scala 169:31]
  assign uart_clock = clock;
  assign uart_reset = reset;
  assign uart_io_rxd = io_rxd; // @[Tile.scala 172:15]
  assign uart_io_rxChannel_ready = uartController_io__rxChannel_ready; // @[Tile.scala 170:31]
  assign uart_io_txChannel_valid = uartController_io__txChannel_valid; // @[Tile.scala 169:31]
  assign uart_io_txChannel_bits = uartController_io__txChannel_bits; // @[Tile.scala 169:31]
  assign rtc_clock = clock;
  assign rtc_reset = reset;
  assign rtc_io_req_valid = regmapper_io_rtc_req_valid; // @[Tile.scala 177:20]
  assign rtc_io_req_bits_addr = regmapper_io_rtc_req_bits_addr; // @[Tile.scala 177:20]
  assign rtc_io_req_bits_data = regmapper_io_rtc_req_bits_data; // @[Tile.scala 177:20]
  assign rtc_io_req_bits_mask = regmapper_io_rtc_req_bits_mask; // @[Tile.scala 177:20]
endmodule
